Sum Block

.include TSMC_180nm.txt
.include gates.cir
.param supply=1.8
.param LAMBDA=0.09u
.param width=10*LAMBDA 
.global gnd vdd

Vrail vdd gnd {supply}
VA A gnd pulse 0 1.8 0ns 100ps 100ps 25ns 50ns
VB B gnd pulse 0 1.8 0ns 100ps 100ps 50ns 100ns
VC C gnd pulse 0 1.8 0ns 100ps 100ps 100ns 200ns

XXOR1 A B p vdd gnd XOR
XXOR2 C p S vdd gnd XOR

.tran 0.1n 200n

.control
run
set color0 = white
set color1 = black
set curplottitle = 'NagamallaSaiAbhinav_2024102037'
plot v(S) v(C)+2 v(B)+4 v(A)+6
.endc