magic
tech scmos
timestamp 1763217344
<< checkpaint >>
rect 227439600 4800 1033480003 23899
rect 227440000 -7 1033480003 4800
<< nwell >>
rect 14 721 48 753
rect -23 644 11 696
rect 55 689 79 721
rect 45 639 81 659
rect 45 607 105 639
rect 112 582 146 614
rect -23 544 11 576
rect -28 470 6 522
rect 45 509 81 561
rect 104 497 162 529
rect 35 451 71 471
rect 35 419 95 451
rect 158 446 194 466
rect -28 370 6 402
rect 109 395 143 427
rect 158 414 218 446
rect -29 297 5 349
rect 26 321 62 373
rect 148 302 206 334
rect 33 260 69 280
rect -29 197 5 229
rect 33 228 93 260
rect 109 203 143 235
rect 153 229 189 249
rect 153 197 213 229
rect -27 97 7 149
rect 33 130 69 182
rect 111 118 169 150
rect 27 72 63 92
rect 169 77 205 97
rect 27 71 87 72
rect 27 40 121 71
rect 169 45 229 77
rect 87 39 121 40
rect -27 -3 7 29
<< ntransistor >>
rect 25 688 27 708
rect 35 688 37 708
rect 66 673 68 683
rect -12 621 -10 631
rect -2 621 0 631
rect -12 590 -10 610
rect -2 590 0 610
rect 57 585 59 595
rect 67 585 69 595
rect 92 589 94 599
rect 123 549 125 569
rect 133 549 135 569
rect 57 487 59 497
rect 67 487 69 497
rect -17 447 -15 457
rect -7 447 -5 457
rect -17 416 -15 436
rect -7 416 -5 436
rect 115 464 117 484
rect 125 464 127 484
rect 149 481 151 491
rect 47 397 49 407
rect 57 397 59 407
rect 82 401 84 411
rect 170 392 172 402
rect 180 392 182 402
rect 205 396 207 406
rect 120 362 122 382
rect 130 362 132 382
rect 38 299 40 309
rect 48 299 50 309
rect -18 274 -16 284
rect -8 274 -6 284
rect -18 243 -16 263
rect -8 243 -6 263
rect 159 269 161 289
rect 169 269 171 289
rect 193 286 195 296
rect 45 206 47 216
rect 55 206 57 216
rect 80 210 82 220
rect 120 170 122 190
rect 130 170 132 190
rect 165 175 167 185
rect 175 175 177 185
rect 200 179 202 189
rect 45 108 47 118
rect 55 108 57 118
rect -16 74 -14 84
rect -6 74 -4 84
rect -16 43 -14 63
rect -6 43 -4 63
rect 122 85 124 105
rect 132 85 134 105
rect 156 102 158 112
rect 39 18 41 28
rect 49 18 51 28
rect 74 22 76 32
rect 98 6 100 26
rect 108 6 110 26
rect 181 23 183 33
rect 191 23 193 33
rect 216 27 218 37
<< ptransistor >>
rect 25 727 27 747
rect 35 727 37 747
rect -12 650 -10 690
rect -2 650 0 690
rect 66 695 68 715
rect 57 613 59 653
rect 67 613 69 653
rect 92 613 94 633
rect 123 588 125 608
rect 133 588 135 608
rect -12 550 -10 570
rect -2 550 0 570
rect -17 476 -15 516
rect -7 476 -5 516
rect 57 515 59 555
rect 67 515 69 555
rect 115 503 117 523
rect 125 503 127 523
rect 149 503 151 523
rect 47 425 49 465
rect 57 425 59 465
rect 82 425 84 445
rect 120 401 122 421
rect 130 401 132 421
rect 170 420 172 460
rect 180 420 182 460
rect 205 420 207 440
rect -17 376 -15 396
rect -7 376 -5 396
rect -18 303 -16 343
rect -8 303 -6 343
rect 38 327 40 367
rect 48 327 50 367
rect 159 308 161 328
rect 169 308 171 328
rect 193 308 195 328
rect 45 234 47 274
rect 55 234 57 274
rect 80 234 82 254
rect -18 203 -16 223
rect -8 203 -6 223
rect 120 209 122 229
rect 130 209 132 229
rect 165 203 167 243
rect 175 203 177 243
rect 200 203 202 223
rect -16 103 -14 143
rect -6 103 -4 143
rect 45 136 47 176
rect 55 136 57 176
rect 122 124 124 144
rect 132 124 134 144
rect 156 124 158 144
rect 39 46 41 86
rect 49 46 51 86
rect 74 46 76 66
rect 98 45 100 65
rect 108 45 110 65
rect 181 51 183 91
rect 191 51 193 91
rect 216 51 218 71
rect -16 3 -14 23
rect -6 3 -4 23
<< ndiffusion >>
rect 20 692 25 708
rect 24 688 25 692
rect 27 688 35 708
rect 37 704 38 708
rect 37 688 42 704
rect 61 677 66 683
rect 65 673 66 677
rect 68 679 69 683
rect 68 673 73 679
rect -17 625 -12 631
rect -13 621 -12 625
rect -10 627 -8 631
rect -4 627 -2 631
rect -10 621 -2 627
rect 0 625 5 631
rect 0 621 1 625
rect -13 606 -12 610
rect -17 590 -12 606
rect -10 590 -2 610
rect 0 594 5 610
rect 0 590 1 594
rect 52 589 57 595
rect 56 585 57 589
rect 59 591 61 595
rect 65 591 67 595
rect 59 585 67 591
rect 69 589 74 595
rect 87 593 92 599
rect 91 589 92 593
rect 94 595 95 599
rect 94 589 99 595
rect 69 585 70 589
rect 118 553 123 569
rect 122 549 123 553
rect 125 549 133 569
rect 135 565 136 569
rect 135 549 140 565
rect 52 491 57 497
rect 56 487 57 491
rect 59 493 61 497
rect 65 493 67 497
rect 59 487 67 493
rect 69 491 74 497
rect 69 487 70 491
rect 144 485 149 491
rect 110 468 115 484
rect -22 451 -17 457
rect -18 447 -17 451
rect -15 453 -13 457
rect -9 453 -7 457
rect -15 447 -7 453
rect -5 451 0 457
rect -5 447 -4 451
rect -18 432 -17 436
rect -22 416 -17 432
rect -15 416 -7 436
rect -5 420 0 436
rect 114 464 115 468
rect 117 464 125 484
rect 127 480 128 484
rect 148 481 149 485
rect 151 487 152 491
rect 151 481 156 487
rect 127 464 132 480
rect -5 416 -4 420
rect 42 401 47 407
rect 46 397 47 401
rect 49 403 51 407
rect 55 403 57 407
rect 49 397 57 403
rect 59 401 64 407
rect 77 405 82 411
rect 81 401 82 405
rect 84 407 85 411
rect 84 401 89 407
rect 59 397 60 401
rect 165 396 170 402
rect 169 392 170 396
rect 172 398 174 402
rect 178 398 180 402
rect 172 392 180 398
rect 182 396 187 402
rect 200 400 205 406
rect 204 396 205 400
rect 207 402 208 406
rect 207 396 212 402
rect 182 392 183 396
rect 115 366 120 382
rect 119 362 120 366
rect 122 362 130 382
rect 132 378 133 382
rect 132 362 137 378
rect 33 303 38 309
rect 37 299 38 303
rect 40 305 42 309
rect 46 305 48 309
rect 40 299 48 305
rect 50 303 55 309
rect 50 299 51 303
rect 188 290 193 296
rect -23 278 -18 284
rect -19 274 -18 278
rect -16 280 -14 284
rect -10 280 -8 284
rect -16 274 -8 280
rect -6 278 -1 284
rect -6 274 -5 278
rect -19 259 -18 263
rect -23 243 -18 259
rect -16 243 -8 263
rect -6 247 -1 263
rect -6 243 -5 247
rect 154 273 159 289
rect 158 269 159 273
rect 161 269 169 289
rect 171 285 172 289
rect 192 286 193 290
rect 195 292 196 296
rect 195 286 200 292
rect 171 269 176 285
rect 40 210 45 216
rect 44 206 45 210
rect 47 212 49 216
rect 53 212 55 216
rect 47 206 55 212
rect 57 210 62 216
rect 75 214 80 220
rect 79 210 80 214
rect 82 216 83 220
rect 82 210 87 216
rect 57 206 58 210
rect 115 174 120 190
rect 119 170 120 174
rect 122 170 130 190
rect 132 186 133 190
rect 132 170 137 186
rect 160 179 165 185
rect 164 175 165 179
rect 167 181 169 185
rect 173 181 175 185
rect 167 175 175 181
rect 177 179 182 185
rect 195 183 200 189
rect 199 179 200 183
rect 202 185 203 189
rect 202 179 207 185
rect 177 175 178 179
rect 40 112 45 118
rect 44 108 45 112
rect 47 114 49 118
rect 53 114 55 118
rect 47 108 55 114
rect 57 112 62 118
rect 57 108 58 112
rect 151 106 156 112
rect 117 89 122 105
rect -21 78 -16 84
rect -17 74 -16 78
rect -14 80 -12 84
rect -8 80 -6 84
rect -14 74 -6 80
rect -4 78 1 84
rect -4 74 -3 78
rect -17 59 -16 63
rect -21 43 -16 59
rect -14 43 -6 63
rect -4 47 1 63
rect -4 43 -3 47
rect 121 85 122 89
rect 124 85 132 105
rect 134 101 135 105
rect 155 102 156 106
rect 158 108 159 112
rect 158 102 163 108
rect 134 85 139 101
rect 34 22 39 28
rect 38 18 39 22
rect 41 24 43 28
rect 47 24 49 28
rect 41 18 49 24
rect 51 22 56 28
rect 69 26 74 32
rect 73 22 74 26
rect 76 28 77 32
rect 76 22 81 28
rect 176 27 181 33
rect 51 18 52 22
rect 93 10 98 26
rect 97 6 98 10
rect 100 6 108 26
rect 110 22 111 26
rect 180 23 181 27
rect 183 29 185 33
rect 189 29 191 33
rect 183 23 191 29
rect 193 27 198 33
rect 211 31 216 37
rect 215 27 216 31
rect 218 33 219 37
rect 218 27 223 33
rect 193 23 194 27
rect 110 6 115 22
<< pdiffusion >>
rect 24 743 25 747
rect 20 727 25 743
rect 27 731 35 747
rect 27 727 29 731
rect 33 727 35 731
rect 37 743 38 747
rect 37 727 42 743
rect 65 711 66 715
rect -13 686 -12 690
rect -17 650 -12 686
rect -10 650 -2 690
rect 0 654 5 690
rect 61 695 66 711
rect 68 699 73 715
rect 68 695 69 699
rect 0 650 1 654
rect 56 649 57 653
rect 52 613 57 649
rect 59 613 67 653
rect 69 617 74 653
rect 69 613 70 617
rect 91 629 92 633
rect 87 613 92 629
rect 94 617 99 633
rect 94 613 95 617
rect 122 604 123 608
rect 118 588 123 604
rect 125 592 133 608
rect 125 588 127 592
rect 131 588 133 592
rect 135 604 136 608
rect 135 588 140 604
rect -17 554 -12 570
rect -13 550 -12 554
rect -10 566 -8 570
rect -4 566 -2 570
rect -10 550 -2 566
rect 0 554 5 570
rect 0 550 1 554
rect 56 551 57 555
rect -18 512 -17 516
rect -22 476 -17 512
rect -15 476 -7 516
rect -5 480 0 516
rect 52 515 57 551
rect 59 515 67 555
rect 69 519 74 555
rect 69 515 70 519
rect 114 519 115 523
rect 110 503 115 519
rect 117 507 125 523
rect 117 503 119 507
rect 123 503 125 507
rect 127 519 128 523
rect 127 503 132 519
rect 148 519 149 523
rect 144 503 149 519
rect 151 507 156 523
rect 151 503 152 507
rect -5 476 -4 480
rect 46 461 47 465
rect 42 425 47 461
rect 49 425 57 465
rect 59 429 64 465
rect 169 456 170 460
rect 59 425 60 429
rect 81 441 82 445
rect 77 425 82 441
rect 84 429 89 445
rect 84 425 85 429
rect 119 417 120 421
rect 115 401 120 417
rect 122 405 130 421
rect 122 401 124 405
rect 128 401 130 405
rect 132 417 133 421
rect 165 420 170 456
rect 172 420 180 460
rect 182 424 187 460
rect 182 420 183 424
rect 204 436 205 440
rect 200 420 205 436
rect 207 424 212 440
rect 207 420 208 424
rect 132 401 137 417
rect -22 380 -17 396
rect -18 376 -17 380
rect -15 392 -13 396
rect -9 392 -7 396
rect -15 376 -7 392
rect -5 380 0 396
rect -5 376 -4 380
rect 37 363 38 367
rect -19 339 -18 343
rect -23 303 -18 339
rect -16 303 -8 343
rect -6 307 -1 343
rect 33 327 38 363
rect 40 327 48 367
rect 50 331 55 367
rect 50 327 51 331
rect 158 324 159 328
rect -6 303 -5 307
rect 154 308 159 324
rect 161 312 169 328
rect 161 308 163 312
rect 167 308 169 312
rect 171 324 172 328
rect 171 308 176 324
rect 192 324 193 328
rect 188 308 193 324
rect 195 312 200 328
rect 195 308 196 312
rect 44 270 45 274
rect 40 234 45 270
rect 47 234 55 274
rect 57 238 62 274
rect 57 234 58 238
rect 79 250 80 254
rect 75 234 80 250
rect 82 238 87 254
rect 82 234 83 238
rect 164 239 165 243
rect -23 207 -18 223
rect -19 203 -18 207
rect -16 219 -14 223
rect -10 219 -8 223
rect -16 203 -8 219
rect -6 207 -1 223
rect 119 225 120 229
rect -6 203 -5 207
rect 115 209 120 225
rect 122 213 130 229
rect 122 209 124 213
rect 128 209 130 213
rect 132 225 133 229
rect 132 209 137 225
rect 160 203 165 239
rect 167 203 175 243
rect 177 207 182 243
rect 177 203 178 207
rect 199 219 200 223
rect 195 203 200 219
rect 202 207 207 223
rect 202 203 203 207
rect 44 172 45 176
rect -17 139 -16 143
rect -21 103 -16 139
rect -14 103 -6 143
rect -4 107 1 143
rect 40 136 45 172
rect 47 136 55 176
rect 57 140 62 176
rect 57 136 58 140
rect 121 140 122 144
rect 117 124 122 140
rect 124 128 132 144
rect 124 124 126 128
rect 130 124 132 128
rect 134 140 135 144
rect 134 124 139 140
rect 155 140 156 144
rect 151 124 156 140
rect 158 128 163 144
rect 158 124 159 128
rect -4 103 -3 107
rect 38 82 39 86
rect 34 46 39 82
rect 41 46 49 86
rect 51 50 56 86
rect 180 87 181 91
rect 51 46 52 50
rect 73 62 74 66
rect 69 46 74 62
rect 76 50 81 66
rect 76 46 77 50
rect 97 61 98 65
rect 93 45 98 61
rect 100 49 108 65
rect 100 45 102 49
rect 106 45 108 49
rect 110 61 111 65
rect 110 45 115 61
rect 176 51 181 87
rect 183 51 191 91
rect 193 55 198 91
rect 193 51 194 55
rect 215 67 216 71
rect 211 51 216 67
rect 218 55 223 71
rect 218 51 219 55
rect -21 7 -16 23
rect -17 3 -16 7
rect -14 19 -12 23
rect -8 19 -6 23
rect -14 3 -6 19
rect -4 7 1 23
rect -4 3 -3 7
<< ndcontact >>
rect 20 688 24 692
rect 38 704 42 708
rect 61 673 65 677
rect 69 679 73 683
rect -17 621 -13 625
rect -8 627 -4 631
rect 1 621 5 625
rect -17 606 -13 610
rect 1 590 5 594
rect 52 585 56 589
rect 61 591 65 595
rect 87 589 91 593
rect 95 595 99 599
rect 70 585 74 589
rect 118 549 122 553
rect 136 565 140 569
rect 52 487 56 491
rect 61 493 65 497
rect 70 487 74 491
rect -22 447 -18 451
rect -13 453 -9 457
rect -4 447 0 451
rect -22 432 -18 436
rect 110 464 114 468
rect 128 480 132 484
rect 144 481 148 485
rect 152 487 156 491
rect -4 416 0 420
rect 42 397 46 401
rect 51 403 55 407
rect 77 401 81 405
rect 85 407 89 411
rect 60 397 64 401
rect 165 392 169 396
rect 174 398 178 402
rect 200 396 204 400
rect 208 402 212 406
rect 183 392 187 396
rect 115 362 119 366
rect 133 378 137 382
rect 33 299 37 303
rect 42 305 46 309
rect 51 299 55 303
rect -23 274 -19 278
rect -14 280 -10 284
rect -5 274 -1 278
rect -23 259 -19 263
rect -5 243 -1 247
rect 154 269 158 273
rect 172 285 176 289
rect 188 286 192 290
rect 196 292 200 296
rect 40 206 44 210
rect 49 212 53 216
rect 75 210 79 214
rect 83 216 87 220
rect 58 206 62 210
rect 115 170 119 174
rect 133 186 137 190
rect 160 175 164 179
rect 169 181 173 185
rect 195 179 199 183
rect 203 185 207 189
rect 178 175 182 179
rect 40 108 44 112
rect 49 114 53 118
rect 58 108 62 112
rect -21 74 -17 78
rect -12 80 -8 84
rect -3 74 1 78
rect -21 59 -17 63
rect -3 43 1 47
rect 117 85 121 89
rect 135 101 139 105
rect 151 102 155 106
rect 159 108 163 112
rect 34 18 38 22
rect 43 24 47 28
rect 69 22 73 26
rect 77 28 81 32
rect 52 18 56 22
rect 93 6 97 10
rect 111 22 115 26
rect 176 23 180 27
rect 185 29 189 33
rect 211 27 215 31
rect 219 33 223 37
rect 194 23 198 27
<< pdcontact >>
rect 20 743 24 747
rect 29 727 33 731
rect 38 743 42 747
rect 61 711 65 715
rect -17 686 -13 690
rect 69 695 73 699
rect 1 650 5 654
rect 52 649 56 653
rect 70 613 74 617
rect 87 629 91 633
rect 95 613 99 617
rect 118 604 122 608
rect 127 588 131 592
rect 136 604 140 608
rect -17 550 -13 554
rect -8 566 -4 570
rect 1 550 5 554
rect 52 551 56 555
rect -22 512 -18 516
rect 70 515 74 519
rect 110 519 114 523
rect 119 503 123 507
rect 128 519 132 523
rect 144 519 148 523
rect 152 503 156 507
rect -4 476 0 480
rect 42 461 46 465
rect 165 456 169 460
rect 60 425 64 429
rect 77 441 81 445
rect 85 425 89 429
rect 115 417 119 421
rect 124 401 128 405
rect 133 417 137 421
rect 183 420 187 424
rect 200 436 204 440
rect 208 420 212 424
rect -22 376 -18 380
rect -13 392 -9 396
rect -4 376 0 380
rect 33 363 37 367
rect -23 339 -19 343
rect 51 327 55 331
rect 154 324 158 328
rect -5 303 -1 307
rect 163 308 167 312
rect 172 324 176 328
rect 188 324 192 328
rect 196 308 200 312
rect 40 270 44 274
rect 58 234 62 238
rect 75 250 79 254
rect 83 234 87 238
rect 160 239 164 243
rect -23 203 -19 207
rect -14 219 -10 223
rect 115 225 119 229
rect -5 203 -1 207
rect 124 209 128 213
rect 133 225 137 229
rect 178 203 182 207
rect 195 219 199 223
rect 203 203 207 207
rect 40 172 44 176
rect -21 139 -17 143
rect 58 136 62 140
rect 117 140 121 144
rect 126 124 130 128
rect 135 140 139 144
rect 151 140 155 144
rect 159 124 163 128
rect -3 103 1 107
rect 34 82 38 86
rect 176 87 180 91
rect 52 46 56 50
rect 69 62 73 66
rect 77 46 81 50
rect 93 61 97 65
rect 102 45 106 49
rect 111 61 115 65
rect 194 51 198 55
rect 211 67 215 71
rect 219 51 223 55
rect -21 3 -17 7
rect -12 19 -8 23
rect -3 3 1 7
<< polysilicon >>
rect 25 747 27 751
rect 35 747 37 751
rect 25 708 27 727
rect 35 708 37 727
rect 66 715 68 718
rect -12 690 -10 693
rect -2 690 0 693
rect 25 685 27 688
rect 35 685 37 688
rect 66 683 68 695
rect 66 670 68 673
rect 57 653 59 656
rect 67 653 69 656
rect -12 631 -10 650
rect -2 631 0 650
rect -12 618 -10 621
rect -2 618 0 621
rect 92 633 94 636
rect -12 610 -10 613
rect -2 610 0 613
rect 57 595 59 613
rect 67 595 69 613
rect 92 599 94 613
rect 123 608 125 612
rect 133 608 135 612
rect -12 570 -10 590
rect -2 570 0 590
rect 92 586 94 589
rect 57 582 59 585
rect 67 582 69 585
rect 123 569 125 588
rect 133 569 135 588
rect 57 555 59 558
rect 67 555 69 558
rect -12 546 -10 550
rect -2 546 0 550
rect -17 516 -15 519
rect -7 516 -5 519
rect 123 546 125 549
rect 133 546 135 549
rect 115 523 117 527
rect 125 523 127 527
rect 149 523 151 526
rect 57 497 59 515
rect 67 497 69 515
rect 57 484 59 487
rect 67 484 69 487
rect 115 484 117 503
rect 125 484 127 503
rect 149 491 151 503
rect -17 457 -15 476
rect -7 457 -5 476
rect 47 465 49 468
rect 57 465 59 468
rect -17 444 -15 447
rect -7 444 -5 447
rect -17 436 -15 439
rect -7 436 -5 439
rect 149 478 151 481
rect 115 461 117 464
rect 125 461 127 464
rect 170 460 172 463
rect 180 460 182 463
rect 82 445 84 448
rect -17 396 -15 416
rect -7 396 -5 416
rect 47 407 49 425
rect 57 407 59 425
rect 82 411 84 425
rect 120 421 122 425
rect 130 421 132 425
rect 205 440 207 443
rect 170 402 172 420
rect 180 402 182 420
rect 205 406 207 420
rect 82 398 84 401
rect 47 394 49 397
rect 57 394 59 397
rect 120 382 122 401
rect 130 382 132 401
rect 205 393 207 396
rect 170 389 172 392
rect 180 389 182 392
rect -17 372 -15 376
rect -7 372 -5 376
rect 38 367 40 370
rect 48 367 50 370
rect -18 343 -16 346
rect -8 343 -6 346
rect 120 359 122 362
rect 130 359 132 362
rect 159 328 161 332
rect 169 328 171 332
rect 193 328 195 331
rect 38 309 40 327
rect 48 309 50 327
rect -18 284 -16 303
rect -8 284 -6 303
rect 38 296 40 299
rect 48 296 50 299
rect 159 289 161 308
rect 169 289 171 308
rect 193 296 195 308
rect 45 274 47 277
rect 55 274 57 277
rect -18 271 -16 274
rect -8 271 -6 274
rect -18 263 -16 266
rect -8 263 -6 266
rect -18 223 -16 243
rect -8 223 -6 243
rect 193 283 195 286
rect 159 266 161 269
rect 169 266 171 269
rect 80 254 82 257
rect 165 243 167 246
rect 175 243 177 246
rect 45 216 47 234
rect 55 216 57 234
rect 80 220 82 234
rect 120 229 122 233
rect 130 229 132 233
rect 80 207 82 210
rect 45 203 47 206
rect 55 203 57 206
rect -18 199 -16 203
rect -8 199 -6 203
rect 120 190 122 209
rect 130 190 132 209
rect 200 223 202 226
rect 45 176 47 179
rect 55 176 57 179
rect -16 143 -14 146
rect -6 143 -4 146
rect 165 185 167 203
rect 175 185 177 203
rect 200 189 202 203
rect 200 176 202 179
rect 165 172 167 175
rect 175 172 177 175
rect 120 167 122 170
rect 130 167 132 170
rect 122 144 124 148
rect 132 144 134 148
rect 156 144 158 147
rect 45 118 47 136
rect 55 118 57 136
rect 45 105 47 108
rect 55 105 57 108
rect 122 105 124 124
rect 132 105 134 124
rect 156 112 158 124
rect -16 84 -14 103
rect -6 84 -4 103
rect 39 86 41 89
rect 49 86 51 89
rect -16 71 -14 74
rect -6 71 -4 74
rect -16 63 -14 66
rect -6 63 -4 66
rect 156 99 158 102
rect 181 91 183 94
rect 191 91 193 94
rect 122 82 124 85
rect 132 82 134 85
rect 74 66 76 69
rect 98 65 100 69
rect 108 65 110 69
rect -16 23 -14 43
rect -6 23 -4 43
rect 39 28 41 46
rect 49 28 51 46
rect 74 32 76 46
rect 216 71 218 74
rect 98 26 100 45
rect 108 26 110 45
rect 181 33 183 51
rect 191 33 193 51
rect 216 37 218 51
rect 74 19 76 22
rect 39 15 41 18
rect 49 15 51 18
rect 216 24 218 27
rect 181 20 183 23
rect 191 20 193 23
rect 98 3 100 6
rect 108 3 110 6
rect -16 -1 -14 3
rect -6 -1 -4 3
<< polycontact >>
rect 21 716 25 720
rect 31 709 35 713
rect 62 684 66 688
rect -16 632 -12 636
rect -6 639 -2 643
rect 53 596 57 600
rect 63 602 67 606
rect 88 600 92 604
rect -16 577 -12 581
rect -6 585 -2 589
rect 119 577 123 581
rect 129 570 133 574
rect 53 498 57 502
rect 63 504 67 508
rect 111 492 115 496
rect 121 485 125 489
rect 145 492 149 496
rect -21 458 -17 462
rect -11 465 -7 469
rect -21 403 -17 407
rect -11 411 -7 415
rect 43 408 47 412
rect 53 414 57 418
rect 78 412 82 416
rect 166 403 170 407
rect 176 409 180 413
rect 201 407 205 411
rect 116 390 120 394
rect 126 383 130 387
rect 34 310 38 314
rect 44 316 48 320
rect -22 285 -18 289
rect -12 292 -8 296
rect 155 297 159 301
rect 165 290 169 294
rect 189 297 193 301
rect -22 230 -18 234
rect -12 238 -8 242
rect 41 217 45 221
rect 51 223 55 227
rect 76 221 80 225
rect 116 198 120 202
rect 126 191 130 195
rect 161 186 165 190
rect 171 192 175 196
rect 196 190 200 194
rect 41 119 45 123
rect 51 125 55 129
rect 118 113 122 117
rect 128 106 132 110
rect 152 113 156 117
rect -20 85 -16 89
rect -10 92 -6 96
rect -20 30 -16 34
rect -10 38 -6 42
rect 35 29 39 33
rect 45 35 49 39
rect 70 33 74 37
rect 94 34 98 38
rect 104 27 108 31
rect 177 34 181 38
rect 187 40 191 44
rect 212 38 216 42
<< metal1 >>
rect 20 754 42 757
rect 20 747 23 754
rect 39 747 42 754
rect 14 716 21 719
rect 30 719 33 727
rect 56 722 66 725
rect 30 716 48 719
rect 14 709 31 712
rect 39 708 42 716
rect -23 696 6 700
rect -17 690 -13 696
rect 20 685 23 688
rect 45 687 48 716
rect 61 715 64 722
rect 70 688 73 695
rect 19 682 24 685
rect 41 684 62 687
rect 70 685 110 688
rect -32 639 -6 643
rect -32 581 -29 639
rect 1 636 5 650
rect -26 632 -16 636
rect -8 632 32 636
rect -26 589 -23 632
rect -8 631 -4 632
rect -17 617 -13 621
rect 1 617 5 621
rect -17 614 5 617
rect -17 610 -13 614
rect 28 599 32 632
rect 45 606 48 684
rect 70 683 73 685
rect 61 669 64 673
rect 61 666 71 669
rect 52 660 85 663
rect 52 653 55 660
rect 82 643 85 660
rect 82 640 90 643
rect 87 633 90 640
rect 45 603 63 606
rect 71 604 74 613
rect 96 604 99 613
rect 118 615 140 618
rect 118 608 121 615
rect 137 608 140 615
rect 71 601 88 604
rect 28 596 38 599
rect 43 596 53 599
rect 71 599 74 601
rect 96 601 105 604
rect 96 599 99 601
rect 62 596 74 599
rect 62 595 65 596
rect -26 585 -6 589
rect 1 581 5 590
rect -32 577 -16 581
rect -8 577 27 581
rect -8 570 -4 577
rect 23 573 27 577
rect 52 579 55 585
rect 71 579 74 585
rect 87 579 90 589
rect 52 576 90 579
rect 102 580 105 601
rect 102 577 119 580
rect 128 580 131 588
rect 128 577 149 580
rect 20 570 129 573
rect 137 569 140 577
rect 50 564 56 567
rect 52 555 55 564
rect -17 542 -13 550
rect 1 544 5 550
rect 118 546 121 549
rect 1 542 6 544
rect -17 539 6 542
rect 117 543 122 546
rect 110 530 147 533
rect -28 522 1 526
rect 110 523 113 530
rect 129 523 132 530
rect -22 516 -18 522
rect 144 523 147 530
rect 44 505 63 508
rect 71 506 74 515
rect 71 503 82 506
rect 8 498 24 501
rect 29 498 53 501
rect 71 501 74 503
rect 62 498 74 501
rect -37 465 -11 469
rect -37 407 -34 465
rect -4 462 0 476
rect 8 462 11 498
rect -31 458 -21 462
rect -13 458 11 462
rect -31 415 -28 458
rect -13 457 -9 458
rect -22 443 -18 447
rect -4 443 0 447
rect -22 440 0 443
rect -22 436 -18 440
rect -31 411 -11 415
rect -4 407 0 416
rect 35 418 38 498
rect 62 497 65 498
rect 52 481 55 487
rect 71 481 74 487
rect 79 488 82 503
rect 100 492 111 495
rect 120 495 123 503
rect 153 496 156 503
rect 120 492 145 495
rect 153 493 162 496
rect 79 485 121 488
rect 129 484 132 492
rect 153 491 156 493
rect 52 478 74 481
rect 42 472 75 475
rect 42 465 45 472
rect 72 455 75 472
rect 110 461 113 464
rect 144 461 147 481
rect 109 458 147 461
rect 72 452 80 455
rect 77 445 80 452
rect 35 415 53 418
rect 61 416 64 425
rect 86 416 89 425
rect 115 428 137 431
rect 115 421 118 428
rect 134 421 137 428
rect 61 413 78 416
rect 22 408 43 411
rect 61 411 64 413
rect 86 413 95 416
rect 159 413 162 493
rect 165 467 198 470
rect 165 460 168 467
rect 195 450 198 467
rect 195 447 203 450
rect 200 440 203 447
rect 86 411 89 413
rect 52 408 64 411
rect 52 407 55 408
rect -37 403 -21 407
rect -13 403 12 407
rect -13 396 -9 403
rect 9 385 12 403
rect 42 391 45 397
rect 61 391 64 397
rect 77 391 80 401
rect 42 388 80 391
rect 92 393 95 413
rect 158 410 176 413
rect 184 411 187 420
rect 209 411 212 420
rect 184 408 201 411
rect 92 390 116 393
rect 125 393 128 401
rect 154 403 166 406
rect 184 406 187 408
rect 209 408 218 411
rect 209 406 212 408
rect 175 403 187 406
rect 154 393 157 403
rect 175 402 178 403
rect 125 390 157 393
rect 9 382 33 385
rect 108 385 126 386
rect 38 383 126 385
rect 38 382 111 383
rect 134 382 137 390
rect 165 386 168 392
rect 184 386 187 392
rect 200 386 203 396
rect 165 383 203 386
rect -22 368 -18 376
rect 31 376 37 379
rect -4 370 0 376
rect -4 368 1 370
rect -22 365 1 368
rect 33 367 36 376
rect 115 359 118 362
rect 114 356 119 359
rect -29 349 0 353
rect -23 343 -19 349
rect 154 335 191 338
rect 25 317 44 320
rect 52 318 55 327
rect 154 328 157 335
rect 173 328 176 335
rect 188 328 191 335
rect 52 315 105 318
rect 8 310 34 313
rect 52 313 55 315
rect 43 310 55 313
rect -38 292 -12 296
rect -38 234 -35 292
rect -5 289 -1 303
rect 8 289 12 310
rect -32 285 -22 289
rect -14 285 12 289
rect -32 242 -29 285
rect -14 284 -10 285
rect -23 270 -19 274
rect -5 270 -1 274
rect -23 267 -1 270
rect -23 263 -19 267
rect -32 238 -12 242
rect -5 234 -1 243
rect -38 230 -22 234
rect -14 230 9 234
rect -14 223 -10 230
rect 21 220 24 310
rect 43 309 46 310
rect 33 293 36 299
rect 52 293 55 299
rect 33 290 55 293
rect 102 293 105 315
rect 146 297 155 300
rect 164 300 167 308
rect 197 301 200 308
rect 164 297 189 300
rect 197 298 206 301
rect 102 290 165 293
rect 173 289 176 297
rect 197 296 200 298
rect 40 281 73 284
rect 40 274 43 281
rect 70 264 73 281
rect 154 266 157 269
rect 188 266 191 286
rect 70 261 78 264
rect 153 263 191 266
rect 75 254 78 261
rect 203 260 206 298
rect 154 257 206 260
rect 32 224 51 227
rect 59 225 62 234
rect 84 225 87 234
rect 115 236 137 239
rect 115 229 118 236
rect 134 229 137 236
rect 59 222 76 225
rect 21 217 41 220
rect 59 220 62 222
rect 84 222 93 225
rect 84 220 87 222
rect 50 217 62 220
rect -23 195 -19 203
rect -5 197 -1 203
rect -5 195 0 197
rect -23 192 0 195
rect -27 149 2 153
rect -21 143 -17 149
rect 21 129 24 217
rect 50 216 53 217
rect 40 200 43 206
rect 59 200 62 206
rect 75 200 78 210
rect 40 197 78 200
rect 90 201 93 222
rect 90 198 116 201
rect 125 201 128 209
rect 125 198 143 201
rect 33 191 126 194
rect 134 190 137 198
rect 38 185 44 188
rect 140 189 143 198
rect 154 196 157 257
rect 160 250 193 253
rect 160 243 163 250
rect 190 233 193 250
rect 190 230 198 233
rect 195 223 198 230
rect 154 193 171 196
rect 179 194 182 203
rect 204 194 207 203
rect 179 191 196 194
rect 140 186 161 189
rect 179 189 182 191
rect 204 191 213 194
rect 204 189 207 191
rect 170 186 182 189
rect 170 185 173 186
rect 40 176 43 185
rect 115 167 118 170
rect 160 169 163 175
rect 179 169 182 175
rect 195 169 198 179
rect 114 164 119 167
rect 160 166 198 169
rect 117 151 154 154
rect 117 144 120 151
rect 136 144 139 151
rect 151 144 154 151
rect 21 126 51 129
rect 59 127 62 136
rect 59 124 94 127
rect 21 119 41 122
rect 59 122 62 124
rect 50 119 62 122
rect -36 92 -10 96
rect -36 34 -33 92
rect -3 89 1 103
rect 21 89 24 119
rect 50 118 53 119
rect 40 102 43 108
rect 59 102 62 108
rect 91 109 94 124
rect 110 113 118 116
rect 127 116 130 124
rect 160 117 163 124
rect 127 113 152 116
rect 160 114 169 117
rect 91 106 128 109
rect 136 105 139 113
rect 160 112 163 114
rect 40 99 62 102
rect -30 85 -20 89
rect -12 85 24 89
rect -30 42 -27 85
rect -12 84 -8 85
rect -21 70 -17 74
rect -3 70 1 74
rect -21 67 1 70
rect -21 63 -17 67
rect 21 55 24 85
rect 34 93 67 96
rect 34 86 37 93
rect 64 76 67 93
rect 117 82 120 85
rect 151 82 154 102
rect 116 79 154 82
rect 64 73 72 76
rect 69 66 72 73
rect 93 72 115 75
rect 93 65 96 72
rect 112 65 115 72
rect 13 52 24 55
rect -30 38 -10 42
rect -3 34 1 43
rect -36 30 -20 34
rect -12 30 7 34
rect -12 23 -8 30
rect -21 -5 -17 3
rect -3 -3 1 3
rect 4 3 7 30
rect 13 32 16 52
rect 25 36 45 39
rect 53 37 56 46
rect 78 37 81 46
rect 53 34 70 37
rect 13 29 35 32
rect 53 32 56 34
rect 78 34 94 37
rect 103 37 106 45
rect 166 44 169 114
rect 176 98 209 101
rect 176 91 179 98
rect 206 81 209 98
rect 206 78 214 81
rect 211 71 214 78
rect 166 41 187 44
rect 195 42 198 51
rect 220 42 223 51
rect 195 39 212 42
rect 103 34 177 37
rect 195 37 198 39
rect 220 39 229 42
rect 220 37 223 39
rect 186 34 198 37
rect 78 32 81 34
rect 44 29 56 32
rect 44 28 47 29
rect 84 27 104 30
rect 34 12 37 18
rect 53 12 56 18
rect 69 12 72 22
rect 34 9 72 12
rect 84 3 87 27
rect 112 26 115 34
rect 186 33 189 34
rect 176 17 179 23
rect 195 17 198 23
rect 211 17 214 27
rect 176 14 214 17
rect 93 3 96 6
rect 4 0 87 3
rect 92 0 97 3
rect -3 -5 2 -3
rect -21 -8 2 -5
<< m2contact >>
rect 6 696 11 701
rect 110 685 115 690
rect 38 594 43 599
rect 149 577 154 582
rect 15 568 20 573
rect 6 539 11 544
rect 1 522 6 527
rect 39 505 44 510
rect 24 498 29 503
rect 17 408 22 413
rect 218 408 223 413
rect 33 382 38 387
rect 1 365 6 370
rect 0 349 5 354
rect 20 317 25 322
rect 9 230 14 235
rect 141 297 146 302
rect 27 224 32 229
rect 0 192 5 197
rect 2 149 7 154
rect 27 191 33 197
rect 105 113 110 118
rect 20 36 25 41
rect 2 -8 7 -3
<< psm12contact >>
rect 95 492 100 497
<< metal2 >>
rect 8 544 11 696
rect 3 370 6 522
rect 17 413 20 568
rect 40 510 43 594
rect 110 507 113 685
rect 95 504 113 507
rect 2 197 5 349
rect 26 327 29 498
rect 95 497 98 504
rect 20 324 29 327
rect 20 322 26 324
rect 35 232 38 382
rect 151 309 154 577
rect 143 306 154 309
rect 143 302 146 306
rect 11 194 14 230
rect 27 229 38 232
rect 11 191 27 194
rect 4 -3 7 149
rect 27 51 30 191
rect 220 160 223 408
rect 105 157 223 160
rect 105 118 108 157
rect 22 48 30 51
rect 22 41 25 48
<< labels >>
rlabel metal1 60 724 60 724 4 vdd
rlabel metal1 67 667 67 667 1 gnd
rlabel metal1 76 686 76 686 7 c1
rlabel metal1 62 577 62 577 1 gnd
rlabel metal1 67 661 67 661 5 vdd
rlabel metal1 42 685 42 685 3 g0_bar
rlabel metal1 29 597 29 597 3 p1_bar
rlabel metal1 129 616 129 616 5 vdd
rlabel metal1 120 544 120 544 1 gnd
rlabel metal1 29 571 29 571 3 g1_bar
rlabel metal1 143 579 143 579 7 c2
rlabel metal1 53 566 53 566 5 vdd
rlabel metal1 62 479 62 479 1 gnd
rlabel metal1 16 499 16 499 3 p2_bar
rlabel metal1 52 389 52 389 1 gnd
rlabel metal1 57 473 57 473 5 vdd
rlabel metal1 125 532 125 532 1 vdd
rlabel metal1 130 459 130 459 1 gnd
rlabel metal1 117 357 117 357 1 gnd
rlabel metal1 126 429 126 429 5 vdd
rlabel metal1 180 469 180 469 1 vdd
rlabel metal1 181 384 181 384 1 gnd
rlabel metal1 33 377 33 377 1 vdd
rlabel metal1 42 291 42 291 1 gnd
rlabel metal1 53 282 53 282 1 vdd
rlabel metal1 58 198 58 198 1 gnd
rlabel metal1 125 237 125 237 1 vdd
rlabel metal1 117 165 117 165 1 gnd
rlabel metal1 215 409 215 409 7 c3
rlabel metal1 169 337 169 337 1 vdd
rlabel metal1 174 265 174 265 1 gnd
rlabel metal1 179 167 179 167 1 gnd
rlabel metal1 177 251 177 251 1 vdd
rlabel metal1 211 192 211 192 1 c4
rlabel metal1 42 192 42 192 1 g3_bar
rlabel metal1 40 186 40 186 1 vdd
rlabel metal1 48 100 48 100 1 gnd
rlabel metal1 22 120 22 120 1 p4_bar
rlabel metal1 49 94 49 94 1 vdd
rlabel metal1 54 10 54 10 1 gnd
rlabel metal1 12 1 12 1 1 g4_bar
rlabel metal1 133 152 133 152 1 vdd
rlabel metal1 135 80 135 80 1 gnd
rlabel metal1 93 1 93 1 1 gnd
rlabel metal1 104 73 104 73 1 vdd
rlabel metal1 196 15 196 15 1 gnd
rlabel metal1 192 99 192 99 1 vdd
rlabel metal1 226 40 226 40 7 c5
rlabel metal1 -7 698 -7 698 5 vdd
rlabel metal1 -6 616 -6 616 1 gnd
rlabel metal1 -25 609 -25 609 1 b1
rlabel metal1 -31 609 -31 609 3 a1
rlabel metal1 31 755 31 755 5 vdd
rlabel metal1 21 683 21 683 1 gnd
rlabel metal1 15 717 15 717 1 a0
rlabel metal1 15 710 15 710 1 b0
rlabel metal1 12 383 12 383 1 g2_bar
rlabel metal1 -12 524 -12 524 1 vdd
rlabel metal1 -11 441 -11 441 1 gnd
rlabel metal1 -30 433 -30 433 1 b2
rlabel metal1 -36 433 -36 433 3 a2
rlabel metal1 17 311 17 311 1 p3_bar
rlabel metal1 -14 351 -14 351 1 vdd
rlabel metal1 -12 268 -12 268 1 gnd
rlabel metal1 -30 266 -30 266 1 b3
rlabel metal1 -37 266 -37 266 3 a3
rlabel metal1 -14 150 -14 150 1 vdd
rlabel metal1 -10 68 -10 68 1 gnd
rlabel metal1 -29 64 -29 64 1 b4
rlabel metal1 -35 64 -35 64 3 a4
<< end >>
