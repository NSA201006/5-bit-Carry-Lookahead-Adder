magic
tech scmos
timestamp 1763534783
<< checkpaint >>
rect 76322400 6000 950160835 22047
rect 76322800 -7 950160835 6000
<< nwell >>
rect -101 831 -36 863
rect -101 811 -71 831
rect -17 827 9 859
rect 216 820 240 852
rect 302 818 367 850
rect 302 798 332 818
rect 386 814 412 846
rect -101 720 -36 752
rect -101 700 -71 720
rect -17 716 9 748
rect 54 729 88 761
rect 206 730 230 762
rect 246 736 270 768
rect -214 660 -149 692
rect -214 640 -184 660
rect -130 656 -104 688
rect 17 652 51 704
rect 95 697 119 729
rect 319 712 343 744
rect 398 718 422 750
rect 85 647 121 667
rect 85 615 145 647
rect 309 622 333 654
rect 349 628 373 660
rect 388 628 412 660
rect 428 634 452 666
rect 460 663 525 695
rect 460 643 490 663
rect 544 659 570 691
rect -111 581 -46 613
rect -111 561 -81 581
rect -27 577 -1 609
rect 152 590 186 622
rect 17 552 51 584
rect -222 519 -157 551
rect -222 499 -192 519
rect -138 515 -112 547
rect 12 478 46 530
rect 85 517 121 569
rect 317 540 341 572
rect 408 540 432 572
rect 144 505 202 537
rect 75 459 111 479
rect -113 420 -48 452
rect -113 400 -83 420
rect -29 416 -3 448
rect 75 427 135 459
rect 198 454 234 474
rect -237 366 -172 398
rect -237 346 -207 366
rect -153 362 -127 394
rect 12 378 46 410
rect 149 403 183 435
rect 198 422 258 454
rect 307 450 331 482
rect 347 456 371 488
rect 398 450 422 482
rect 438 456 462 488
rect 472 485 537 517
rect 472 465 502 485
rect 556 481 582 513
rect 11 305 45 357
rect 66 329 102 381
rect 322 374 346 406
rect 409 374 433 406
rect 188 310 246 342
rect 472 328 537 360
rect -120 247 -55 279
rect -120 227 -90 247
rect -36 243 -10 275
rect 73 268 109 288
rect 312 284 336 316
rect 352 290 376 322
rect 399 284 423 316
rect 439 290 463 322
rect 472 308 502 328
rect 556 324 582 356
rect 11 205 45 237
rect 73 236 133 268
rect 149 211 183 243
rect 193 237 229 257
rect 193 205 253 237
rect 406 211 430 243
rect 472 209 537 241
rect -238 136 -173 168
rect -238 116 -208 136
rect -154 132 -128 164
rect 13 105 47 157
rect 73 138 109 190
rect 324 169 348 201
rect 472 189 502 209
rect 556 205 582 237
rect 151 126 209 158
rect 396 121 420 153
rect 436 127 460 159
rect -123 49 -58 81
rect 67 80 103 100
rect 209 85 245 105
rect 67 79 127 80
rect -123 29 -93 49
rect -39 45 -13 77
rect 67 48 161 79
rect 209 53 269 85
rect 314 79 338 111
rect 354 85 378 117
rect 475 86 540 118
rect 475 66 505 86
rect 559 82 585 114
rect 127 47 161 48
rect 13 5 47 37
<< ntransistor >>
rect -90 795 -88 805
rect -58 781 -56 821
rect -52 781 -50 821
rect -34 801 -32 821
rect -25 801 -23 821
rect -6 809 -4 819
rect 227 804 229 814
rect 213 772 215 792
rect 242 775 244 795
rect 313 782 315 792
rect 345 768 347 808
rect 351 768 353 808
rect 369 788 371 808
rect 378 788 380 808
rect 397 796 399 806
rect -90 684 -88 694
rect -58 670 -56 710
rect -52 670 -50 710
rect -34 690 -32 710
rect -25 690 -23 710
rect -6 698 -4 708
rect 65 696 67 716
rect 75 696 77 716
rect 217 714 219 724
rect 257 710 259 730
rect 330 696 332 706
rect 409 702 411 712
rect 106 681 108 691
rect 316 664 318 684
rect 345 667 347 687
rect 395 670 397 690
rect 424 673 426 693
rect -203 624 -201 634
rect -171 610 -169 650
rect -165 610 -163 650
rect -147 630 -145 650
rect -138 630 -136 650
rect -119 638 -117 648
rect 28 629 30 639
rect 38 629 40 639
rect 28 598 30 618
rect 38 598 40 618
rect 97 593 99 603
rect 107 593 109 603
rect 132 597 134 607
rect 320 606 322 616
rect 360 602 362 622
rect 399 612 401 622
rect 439 608 441 628
rect 471 627 473 637
rect 503 613 505 653
rect 509 613 511 653
rect 527 633 529 653
rect 536 633 538 653
rect 555 641 557 651
rect -100 545 -98 555
rect -68 531 -66 571
rect -62 531 -60 571
rect -44 551 -42 571
rect -35 551 -33 571
rect -16 559 -14 569
rect -211 483 -209 493
rect -179 469 -177 509
rect -173 469 -171 509
rect -155 489 -153 509
rect -146 489 -144 509
rect -127 497 -125 507
rect 163 557 165 577
rect 173 557 175 577
rect 328 524 330 534
rect 419 524 421 534
rect 97 495 99 505
rect 107 495 109 505
rect 23 455 25 465
rect 33 455 35 465
rect 23 424 25 444
rect 33 424 35 444
rect 155 472 157 492
rect 165 472 167 492
rect 189 489 191 499
rect 314 492 316 512
rect 343 495 345 515
rect 405 492 407 512
rect 434 495 436 515
rect -102 384 -100 394
rect -70 370 -68 410
rect -64 370 -62 410
rect -46 390 -44 410
rect -37 390 -35 410
rect -18 398 -16 408
rect 87 405 89 415
rect 97 405 99 415
rect 122 409 124 419
rect 318 434 320 444
rect 358 430 360 450
rect 409 434 411 444
rect 449 430 451 450
rect 483 449 485 459
rect 515 435 517 475
rect 521 435 523 475
rect 539 455 541 475
rect 548 455 550 475
rect 567 463 569 473
rect 210 400 212 410
rect 220 400 222 410
rect 245 404 247 414
rect -226 330 -224 340
rect -194 316 -192 356
rect -188 316 -186 356
rect -170 336 -168 356
rect -161 336 -159 356
rect -142 344 -140 354
rect 160 370 162 390
rect 170 370 172 390
rect 333 358 335 368
rect 420 358 422 368
rect 78 307 80 317
rect 88 307 90 317
rect 319 326 321 346
rect 348 329 350 349
rect 406 326 408 346
rect 435 329 437 349
rect 22 282 24 292
rect 32 282 34 292
rect 22 251 24 271
rect 32 251 34 271
rect -109 211 -107 221
rect -77 197 -75 237
rect -71 197 -69 237
rect -53 217 -51 237
rect -44 217 -42 237
rect -25 225 -23 235
rect 199 277 201 297
rect 209 277 211 297
rect 233 294 235 304
rect 323 268 325 278
rect 363 264 365 284
rect 483 292 485 302
rect 410 268 412 278
rect 450 264 452 284
rect 515 278 517 318
rect 521 278 523 318
rect 539 298 541 318
rect 548 298 550 318
rect 567 306 569 316
rect 85 214 87 224
rect 95 214 97 224
rect 120 218 122 228
rect -227 100 -225 110
rect -195 86 -193 126
rect -189 86 -187 126
rect -171 106 -169 126
rect -162 106 -160 126
rect -143 114 -141 124
rect 160 178 162 198
rect 170 178 172 198
rect 205 183 207 193
rect 215 183 217 193
rect 240 187 242 197
rect 417 195 419 205
rect 403 163 405 183
rect 432 166 434 186
rect 483 173 485 183
rect 335 153 337 163
rect 515 159 517 199
rect 521 159 523 199
rect 539 179 541 199
rect 548 179 550 199
rect 567 187 569 197
rect 85 116 87 126
rect 95 116 97 126
rect 321 121 323 141
rect 350 124 352 144
rect 24 82 26 92
rect 34 82 36 92
rect 24 51 26 71
rect 34 51 36 71
rect 162 93 164 113
rect 172 93 174 113
rect 196 110 198 120
rect -112 13 -110 23
rect -80 -1 -78 39
rect -74 -1 -72 39
rect -56 19 -54 39
rect -47 19 -45 39
rect -28 27 -26 37
rect 407 105 409 115
rect 447 101 449 121
rect 325 63 327 73
rect 365 59 367 79
rect 79 26 81 36
rect 89 26 91 36
rect 114 30 116 40
rect 486 50 488 60
rect 138 14 140 34
rect 148 14 150 34
rect 221 31 223 41
rect 231 31 233 41
rect 256 35 258 45
rect 518 36 520 76
rect 524 36 526 76
rect 542 56 544 76
rect 551 56 553 76
rect 570 64 572 74
<< ptransistor >>
rect -90 817 -88 857
rect -84 817 -82 857
rect -68 837 -66 857
rect -52 837 -50 857
rect -6 833 -4 853
rect 227 826 229 846
rect 313 804 315 844
rect 319 804 321 844
rect 335 824 337 844
rect 351 824 353 844
rect 397 820 399 840
rect -90 706 -88 746
rect -84 706 -82 746
rect -68 726 -66 746
rect -52 726 -50 746
rect -6 722 -4 742
rect 65 735 67 755
rect 75 735 77 755
rect 217 736 219 756
rect 257 742 259 762
rect -203 646 -201 686
rect -197 646 -195 686
rect -181 666 -179 686
rect -165 666 -163 686
rect -119 662 -117 682
rect 28 658 30 698
rect 38 658 40 698
rect 106 703 108 723
rect 330 718 332 738
rect 409 724 411 744
rect 97 621 99 661
rect 107 621 109 661
rect 132 621 134 641
rect 320 628 322 648
rect 360 634 362 654
rect 399 634 401 654
rect 439 640 441 660
rect 471 649 473 689
rect 477 649 479 689
rect 493 669 495 689
rect 509 669 511 689
rect 555 665 557 685
rect -100 567 -98 607
rect -94 567 -92 607
rect -78 587 -76 607
rect -62 587 -60 607
rect -16 583 -14 603
rect 163 596 165 616
rect 173 596 175 616
rect -211 505 -209 545
rect -205 505 -203 545
rect -189 525 -187 545
rect -173 525 -171 545
rect -127 521 -125 541
rect 28 558 30 578
rect 38 558 40 578
rect 23 484 25 524
rect 33 484 35 524
rect 97 523 99 563
rect 107 523 109 563
rect 328 546 330 566
rect 419 546 421 566
rect 155 511 157 531
rect 165 511 167 531
rect 189 511 191 531
rect -102 406 -100 446
rect -96 406 -94 446
rect -80 426 -78 446
rect -64 426 -62 446
rect -18 422 -16 442
rect 87 433 89 473
rect 97 433 99 473
rect 122 433 124 453
rect -226 352 -224 392
rect -220 352 -218 392
rect -204 372 -202 392
rect -188 372 -186 392
rect -142 368 -140 388
rect 160 409 162 429
rect 170 409 172 429
rect 210 428 212 468
rect 220 428 222 468
rect 318 456 320 476
rect 358 462 360 482
rect 245 428 247 448
rect 409 456 411 476
rect 449 462 451 482
rect 483 471 485 511
rect 489 471 491 511
rect 505 491 507 511
rect 521 491 523 511
rect 567 487 569 507
rect 23 384 25 404
rect 33 384 35 404
rect 22 311 24 351
rect 32 311 34 351
rect 78 335 80 375
rect 88 335 90 375
rect 333 380 335 400
rect 420 380 422 400
rect 199 316 201 336
rect 209 316 211 336
rect 233 316 235 336
rect -109 233 -107 273
rect -103 233 -101 273
rect -87 253 -85 273
rect -71 253 -69 273
rect -25 249 -23 269
rect 85 242 87 282
rect 95 242 97 282
rect 323 290 325 310
rect 363 296 365 316
rect 410 290 412 310
rect 450 296 452 316
rect 483 314 485 354
rect 489 314 491 354
rect 505 334 507 354
rect 521 334 523 354
rect 567 330 569 350
rect 120 242 122 262
rect 22 211 24 231
rect 32 211 34 231
rect 160 217 162 237
rect 170 217 172 237
rect 205 211 207 251
rect 215 211 217 251
rect 240 211 242 231
rect 417 217 419 237
rect -227 122 -225 162
rect -221 122 -219 162
rect -205 142 -203 162
rect -189 142 -187 162
rect -143 138 -141 158
rect 24 111 26 151
rect 34 111 36 151
rect 85 144 87 184
rect 95 144 97 184
rect 483 195 485 235
rect 489 195 491 235
rect 505 215 507 235
rect 521 215 523 235
rect 567 211 569 231
rect 335 175 337 195
rect 162 132 164 152
rect 172 132 174 152
rect 196 132 198 152
rect 407 127 409 147
rect 447 133 449 153
rect -112 35 -110 75
rect -106 35 -104 75
rect -90 55 -88 75
rect -74 55 -72 75
rect -28 51 -26 71
rect 79 54 81 94
rect 89 54 91 94
rect 114 54 116 74
rect 138 53 140 73
rect 148 53 150 73
rect 221 59 223 99
rect 231 59 233 99
rect 325 85 327 105
rect 365 91 367 111
rect 256 59 258 79
rect 486 72 488 112
rect 492 72 494 112
rect 508 92 510 112
rect 524 92 526 112
rect 570 88 572 108
rect 24 11 26 31
rect 34 11 36 31
<< ndiffusion >>
rect -59 817 -58 821
rect -95 799 -90 805
rect -91 795 -90 799
rect -88 801 -87 805
rect -88 795 -83 801
rect -63 781 -58 817
rect -56 781 -52 821
rect -50 785 -45 821
rect -37 817 -34 821
rect -41 801 -34 817
rect -32 801 -25 821
rect -23 805 -15 821
rect -11 813 -6 819
rect -7 809 -6 813
rect -4 815 -1 819
rect -4 809 3 815
rect 222 808 227 814
rect -23 801 -19 805
rect 226 804 227 808
rect 229 810 230 814
rect 229 804 234 810
rect 344 804 345 808
rect -50 781 -49 785
rect 207 777 213 792
rect 212 772 213 777
rect 215 776 220 792
rect 215 772 216 776
rect 236 780 242 795
rect 241 775 242 780
rect 244 779 249 795
rect 308 786 313 792
rect 312 782 313 786
rect 315 788 316 792
rect 315 782 320 788
rect 244 775 245 779
rect 340 768 345 804
rect 347 768 351 808
rect 353 772 358 808
rect 366 804 369 808
rect 362 788 369 804
rect 371 788 378 808
rect 380 792 388 808
rect 392 800 397 806
rect 396 796 397 800
rect 399 802 402 806
rect 399 796 406 802
rect 380 788 384 792
rect 353 768 354 772
rect -59 706 -58 710
rect -95 688 -90 694
rect -91 684 -90 688
rect -88 690 -87 694
rect -88 684 -83 690
rect -63 670 -58 706
rect -56 670 -52 710
rect -50 674 -45 710
rect -37 706 -34 710
rect -41 690 -34 706
rect -32 690 -25 710
rect -23 694 -15 710
rect -11 702 -6 708
rect -7 698 -6 702
rect -4 704 -1 708
rect -4 698 3 704
rect 60 700 65 716
rect -23 690 -19 694
rect -50 670 -49 674
rect 64 696 65 700
rect 67 696 75 716
rect 77 712 78 716
rect 77 696 82 712
rect 212 718 217 724
rect 216 714 217 718
rect 219 720 220 724
rect 219 714 224 720
rect 252 714 257 730
rect 256 710 257 714
rect 259 726 260 730
rect 259 710 264 726
rect 404 706 409 712
rect 325 700 330 706
rect 329 696 330 700
rect 332 702 333 706
rect 408 702 409 706
rect 411 708 412 712
rect 411 702 416 708
rect 332 696 337 702
rect 101 685 106 691
rect 105 681 106 685
rect 108 687 109 691
rect 108 681 113 687
rect 310 669 316 684
rect 315 664 316 669
rect 318 668 323 684
rect 318 664 319 668
rect 339 672 345 687
rect 344 667 345 672
rect 347 671 352 687
rect 347 667 348 671
rect 389 675 395 690
rect 394 670 395 675
rect 397 674 402 690
rect 397 670 398 674
rect 418 678 424 693
rect 423 673 424 678
rect 426 677 431 693
rect 426 673 427 677
rect -172 646 -171 650
rect -208 628 -203 634
rect -204 624 -203 628
rect -201 630 -200 634
rect -201 624 -196 630
rect -176 610 -171 646
rect -169 610 -165 650
rect -163 614 -158 650
rect -150 646 -147 650
rect -154 630 -147 646
rect -145 630 -138 650
rect -136 634 -128 650
rect -124 642 -119 648
rect -120 638 -119 642
rect -117 644 -114 648
rect -117 638 -110 644
rect -136 630 -132 634
rect 23 633 28 639
rect 27 629 28 633
rect 30 635 32 639
rect 36 635 38 639
rect 30 629 38 635
rect 40 633 45 639
rect 40 629 41 633
rect 502 649 503 653
rect -163 610 -162 614
rect 27 614 28 618
rect 23 598 28 614
rect 30 598 38 618
rect 40 602 45 618
rect 466 631 471 637
rect 40 598 41 602
rect 92 597 97 603
rect 96 593 97 597
rect 99 599 101 603
rect 105 599 107 603
rect 99 593 107 599
rect 109 597 114 603
rect 127 601 132 607
rect 131 597 132 601
rect 134 603 135 607
rect 134 597 139 603
rect 109 593 110 597
rect 315 610 320 616
rect 319 606 320 610
rect 322 612 323 616
rect 322 606 327 612
rect 355 606 360 622
rect 359 602 360 606
rect 362 618 363 622
rect 362 602 367 618
rect 394 616 399 622
rect 398 612 399 616
rect 401 618 402 622
rect 401 612 406 618
rect 434 612 439 628
rect 438 608 439 612
rect 441 624 442 628
rect 470 627 471 631
rect 473 633 474 637
rect 473 627 478 633
rect 441 608 446 624
rect 498 613 503 649
rect 505 613 509 653
rect 511 617 516 653
rect 524 649 527 653
rect 520 633 527 649
rect 529 633 536 653
rect 538 637 546 653
rect 550 645 555 651
rect 554 641 555 645
rect 557 647 560 651
rect 557 641 564 647
rect 538 633 542 637
rect 511 613 512 617
rect -69 567 -68 571
rect -105 549 -100 555
rect -101 545 -100 549
rect -98 551 -97 555
rect -98 545 -93 551
rect -73 531 -68 567
rect -66 531 -62 571
rect -60 535 -55 571
rect -47 567 -44 571
rect -51 551 -44 567
rect -42 551 -35 571
rect -33 555 -25 571
rect -21 563 -16 569
rect -17 559 -16 563
rect -14 565 -11 569
rect -14 559 -7 565
rect -33 551 -29 555
rect -60 531 -59 535
rect -180 505 -179 509
rect -216 487 -211 493
rect -212 483 -211 487
rect -209 489 -208 493
rect -209 483 -204 489
rect -184 469 -179 505
rect -177 469 -173 509
rect -171 473 -166 509
rect -158 505 -155 509
rect -162 489 -155 505
rect -153 489 -146 509
rect -144 493 -136 509
rect -132 501 -127 507
rect -128 497 -127 501
rect -125 503 -122 507
rect -125 497 -118 503
rect -144 489 -140 493
rect 158 561 163 577
rect 162 557 163 561
rect 165 557 173 577
rect 175 573 176 577
rect 175 557 180 573
rect 323 528 328 534
rect 327 524 328 528
rect 330 530 331 534
rect 330 524 335 530
rect 414 528 419 534
rect 418 524 419 528
rect 421 530 422 534
rect 421 524 426 530
rect 92 499 97 505
rect 96 495 97 499
rect 99 501 101 505
rect 105 501 107 505
rect 99 495 107 501
rect 109 499 114 505
rect 109 495 110 499
rect 184 493 189 499
rect -171 469 -170 473
rect 150 476 155 492
rect 18 459 23 465
rect 22 455 23 459
rect 25 461 27 465
rect 31 461 33 465
rect 25 455 33 461
rect 35 459 40 465
rect 35 455 36 459
rect 22 440 23 444
rect 18 424 23 440
rect 25 424 33 444
rect 35 428 40 444
rect 154 472 155 476
rect 157 472 165 492
rect 167 488 168 492
rect 188 489 189 493
rect 191 495 192 499
rect 191 489 196 495
rect 308 497 314 512
rect 313 492 314 497
rect 316 496 321 512
rect 316 492 317 496
rect 337 500 343 515
rect 342 495 343 500
rect 345 499 350 515
rect 345 495 346 499
rect 399 497 405 512
rect 404 492 405 497
rect 407 496 412 512
rect 407 492 408 496
rect 428 500 434 515
rect 433 495 434 500
rect 436 499 441 515
rect 436 495 437 499
rect 167 472 172 488
rect 35 424 36 428
rect -71 406 -70 410
rect -107 388 -102 394
rect -103 384 -102 388
rect -100 390 -99 394
rect -100 384 -95 390
rect -75 370 -70 406
rect -68 370 -64 410
rect -62 374 -57 410
rect -49 406 -46 410
rect -53 390 -46 406
rect -44 390 -37 410
rect -35 394 -27 410
rect -23 402 -18 408
rect -19 398 -18 402
rect -16 404 -13 408
rect 82 409 87 415
rect 86 405 87 409
rect 89 411 91 415
rect 95 411 97 415
rect 89 405 97 411
rect 99 409 104 415
rect 117 413 122 419
rect 121 409 122 413
rect 124 415 125 419
rect 124 409 129 415
rect 514 471 515 475
rect 313 438 318 444
rect 317 434 318 438
rect 320 440 321 444
rect 320 434 325 440
rect 353 434 358 450
rect 357 430 358 434
rect 360 446 361 450
rect 360 430 365 446
rect 478 453 483 459
rect 404 438 409 444
rect 408 434 409 438
rect 411 440 412 444
rect 411 434 416 440
rect 444 434 449 450
rect 448 430 449 434
rect 451 446 452 450
rect 482 449 483 453
rect 485 455 486 459
rect 485 449 490 455
rect 451 430 456 446
rect 510 435 515 471
rect 517 435 521 475
rect 523 439 528 475
rect 536 471 539 475
rect 532 455 539 471
rect 541 455 548 475
rect 550 459 558 475
rect 562 467 567 473
rect 566 463 567 467
rect 569 469 572 473
rect 569 463 576 469
rect 550 455 554 459
rect 523 435 524 439
rect 99 405 100 409
rect -16 398 -9 404
rect -35 390 -31 394
rect 205 404 210 410
rect 209 400 210 404
rect 212 406 214 410
rect 218 406 220 410
rect 212 400 220 406
rect 222 404 227 410
rect 240 408 245 414
rect 244 404 245 408
rect 247 410 248 414
rect 247 404 252 410
rect 222 400 223 404
rect -62 370 -61 374
rect -195 352 -194 356
rect -231 334 -226 340
rect -227 330 -226 334
rect -224 336 -223 340
rect -224 330 -219 336
rect -199 316 -194 352
rect -192 316 -188 356
rect -186 320 -181 356
rect -173 352 -170 356
rect -177 336 -170 352
rect -168 336 -161 356
rect -159 340 -151 356
rect -147 348 -142 354
rect -143 344 -142 348
rect -140 350 -137 354
rect -140 344 -133 350
rect -159 336 -155 340
rect -186 316 -185 320
rect 155 374 160 390
rect 159 370 160 374
rect 162 370 170 390
rect 172 386 173 390
rect 172 370 177 386
rect 328 362 333 368
rect 332 358 333 362
rect 335 364 336 368
rect 335 358 340 364
rect 415 362 420 368
rect 419 358 420 362
rect 422 364 423 368
rect 422 358 427 364
rect 73 311 78 317
rect 77 307 78 311
rect 80 313 82 317
rect 86 313 88 317
rect 80 307 88 313
rect 90 311 95 317
rect 313 331 319 346
rect 318 326 319 331
rect 321 330 326 346
rect 321 326 322 330
rect 342 334 348 349
rect 347 329 348 334
rect 350 333 355 349
rect 350 329 351 333
rect 400 331 406 346
rect 405 326 406 331
rect 408 330 413 346
rect 408 326 409 330
rect 429 334 435 349
rect 434 329 435 334
rect 437 333 442 349
rect 437 329 438 333
rect 90 307 91 311
rect 228 298 233 304
rect 17 286 22 292
rect 21 282 22 286
rect 24 288 26 292
rect 30 288 32 292
rect 24 282 32 288
rect 34 286 39 292
rect 34 282 35 286
rect 21 267 22 271
rect 17 251 22 267
rect 24 251 32 271
rect 34 255 39 271
rect 34 251 35 255
rect -78 233 -77 237
rect -114 215 -109 221
rect -110 211 -109 215
rect -107 217 -106 221
rect -107 211 -102 217
rect -82 197 -77 233
rect -75 197 -71 237
rect -69 201 -64 237
rect -56 233 -53 237
rect -60 217 -53 233
rect -51 217 -44 237
rect -42 221 -34 237
rect -30 229 -25 235
rect -26 225 -25 229
rect -23 231 -20 235
rect 194 281 199 297
rect 198 277 199 281
rect 201 277 209 297
rect 211 293 212 297
rect 232 294 233 298
rect 235 300 236 304
rect 235 294 240 300
rect 211 277 216 293
rect 514 314 515 318
rect 478 296 483 302
rect 318 272 323 278
rect 322 268 323 272
rect 325 274 326 278
rect 325 268 330 274
rect 358 268 363 284
rect 362 264 363 268
rect 365 280 366 284
rect 365 264 370 280
rect 482 292 483 296
rect 485 298 486 302
rect 485 292 490 298
rect 405 272 410 278
rect 409 268 410 272
rect 412 274 413 278
rect 412 268 417 274
rect 445 268 450 284
rect 449 264 450 268
rect 452 280 453 284
rect 452 264 457 280
rect 510 278 515 314
rect 517 278 521 318
rect 523 282 528 318
rect 536 314 539 318
rect 532 298 539 314
rect 541 298 548 318
rect 550 302 558 318
rect 562 310 567 316
rect 566 306 567 310
rect 569 312 572 316
rect 569 306 576 312
rect 550 298 554 302
rect 523 278 524 282
rect -23 225 -16 231
rect -42 217 -38 221
rect 80 218 85 224
rect 84 214 85 218
rect 87 220 89 224
rect 93 220 95 224
rect 87 214 95 220
rect 97 218 102 224
rect 115 222 120 228
rect 119 218 120 222
rect 122 224 123 228
rect 122 218 127 224
rect 97 214 98 218
rect -69 197 -68 201
rect -196 122 -195 126
rect -232 104 -227 110
rect -228 100 -227 104
rect -225 106 -224 110
rect -225 100 -220 106
rect -200 86 -195 122
rect -193 86 -189 126
rect -187 90 -182 126
rect -174 122 -171 126
rect -178 106 -171 122
rect -169 106 -162 126
rect -160 110 -152 126
rect -148 118 -143 124
rect -144 114 -143 118
rect -141 120 -138 124
rect -141 114 -134 120
rect 155 182 160 198
rect 159 178 160 182
rect 162 178 170 198
rect 172 194 173 198
rect 172 178 177 194
rect 412 199 417 205
rect 200 187 205 193
rect 204 183 205 187
rect 207 189 209 193
rect 213 189 215 193
rect 207 183 215 189
rect 217 187 222 193
rect 235 191 240 197
rect 239 187 240 191
rect 242 193 243 197
rect 416 195 417 199
rect 419 201 420 205
rect 419 195 424 201
rect 514 195 515 199
rect 242 187 247 193
rect 217 183 218 187
rect 397 168 403 183
rect 402 163 403 168
rect 405 167 410 183
rect 405 163 406 167
rect 426 171 432 186
rect 431 166 432 171
rect 434 170 439 186
rect 478 177 483 183
rect 482 173 483 177
rect 485 179 486 183
rect 485 173 490 179
rect 434 166 435 170
rect 330 157 335 163
rect 334 153 335 157
rect 337 159 338 163
rect 510 159 515 195
rect 517 159 521 199
rect 523 163 528 199
rect 536 195 539 199
rect 532 179 539 195
rect 541 179 548 199
rect 550 183 558 199
rect 562 191 567 197
rect 566 187 567 191
rect 569 193 572 197
rect 569 187 576 193
rect 550 179 554 183
rect 523 159 524 163
rect 337 153 342 159
rect 80 120 85 126
rect 84 116 85 120
rect 87 122 89 126
rect 93 122 95 126
rect 87 116 95 122
rect 97 120 102 126
rect 97 116 98 120
rect 315 126 321 141
rect 320 121 321 126
rect 323 125 328 141
rect 323 121 324 125
rect 344 129 350 144
rect 349 124 350 129
rect 352 128 357 144
rect 352 124 353 128
rect 191 114 196 120
rect -160 106 -156 110
rect 157 97 162 113
rect -187 86 -186 90
rect 19 86 24 92
rect 23 82 24 86
rect 26 88 28 92
rect 32 88 34 92
rect 26 82 34 88
rect 36 86 41 92
rect 36 82 37 86
rect 23 67 24 71
rect 19 51 24 67
rect 26 51 34 71
rect 36 55 41 71
rect 36 51 37 55
rect 161 93 162 97
rect 164 93 172 113
rect 174 109 175 113
rect 195 110 196 114
rect 198 116 199 120
rect 198 110 203 116
rect 174 93 179 109
rect -81 35 -80 39
rect -117 17 -112 23
rect -113 13 -112 17
rect -110 19 -109 23
rect -110 13 -105 19
rect -85 -1 -80 35
rect -78 -1 -74 39
rect -72 3 -67 39
rect -59 35 -56 39
rect -63 19 -56 35
rect -54 19 -47 39
rect -45 23 -37 39
rect -33 31 -28 37
rect -29 27 -28 31
rect -26 33 -23 37
rect -26 27 -19 33
rect 402 109 407 115
rect 406 105 407 109
rect 409 111 410 115
rect 409 105 414 111
rect 442 105 447 121
rect 446 101 447 105
rect 449 117 450 121
rect 449 101 454 117
rect 320 67 325 73
rect 324 63 325 67
rect 327 69 328 73
rect 327 63 332 69
rect 360 63 365 79
rect 364 59 365 63
rect 367 75 368 79
rect 367 59 372 75
rect 517 72 518 76
rect -45 19 -41 23
rect 74 30 79 36
rect 78 26 79 30
rect 81 32 83 36
rect 87 32 89 36
rect 81 26 89 32
rect 91 30 96 36
rect 109 34 114 40
rect 113 30 114 34
rect 116 36 117 40
rect 116 30 121 36
rect 481 54 486 60
rect 485 50 486 54
rect 488 56 489 60
rect 488 50 493 56
rect 216 35 221 41
rect 91 26 92 30
rect 133 18 138 34
rect 137 14 138 18
rect 140 14 148 34
rect 150 30 151 34
rect 220 31 221 35
rect 223 37 225 41
rect 229 37 231 41
rect 223 31 231 37
rect 233 35 238 41
rect 251 39 256 45
rect 255 35 256 39
rect 258 41 259 45
rect 258 35 263 41
rect 513 36 518 72
rect 520 36 524 76
rect 526 40 531 76
rect 539 72 542 76
rect 535 56 542 72
rect 544 56 551 76
rect 553 60 561 76
rect 565 68 570 74
rect 569 64 570 68
rect 572 70 575 74
rect 572 64 579 70
rect 553 56 557 60
rect 526 36 527 40
rect 233 31 234 35
rect 150 14 155 30
rect -72 -1 -71 3
<< pdiffusion >>
rect -91 853 -90 857
rect -95 817 -90 853
rect -88 817 -84 857
rect -82 821 -77 857
rect -69 853 -68 857
rect -73 837 -68 853
rect -66 841 -61 857
rect -66 837 -65 841
rect -53 853 -52 857
rect -57 837 -52 853
rect -50 841 -45 857
rect -50 837 -49 841
rect -7 849 -6 853
rect -11 833 -6 849
rect -4 837 3 853
rect -4 833 -1 837
rect 226 842 227 846
rect 222 826 227 842
rect 229 830 234 846
rect 229 826 230 830
rect 312 840 313 844
rect -82 817 -81 821
rect 308 804 313 840
rect 315 804 319 844
rect 321 808 326 844
rect 334 840 335 844
rect 330 824 335 840
rect 337 828 342 844
rect 337 824 338 828
rect 350 840 351 844
rect 346 824 351 840
rect 353 828 358 844
rect 353 824 354 828
rect 396 836 397 840
rect 392 820 397 836
rect 399 824 406 840
rect 399 820 402 824
rect 321 804 322 808
rect 256 758 257 762
rect 64 751 65 755
rect -91 742 -90 746
rect -95 706 -90 742
rect -88 706 -84 746
rect -82 710 -77 746
rect -69 742 -68 746
rect -73 726 -68 742
rect -66 730 -61 746
rect -66 726 -65 730
rect -53 742 -52 746
rect -57 726 -52 742
rect -50 730 -45 746
rect -50 726 -49 730
rect -7 738 -6 742
rect -11 722 -6 738
rect -4 726 3 742
rect 60 735 65 751
rect 67 739 75 755
rect 67 735 69 739
rect 73 735 75 739
rect 77 751 78 755
rect 77 735 82 751
rect 216 752 217 756
rect 212 736 217 752
rect 219 740 224 756
rect 252 742 257 758
rect 259 746 264 762
rect 259 742 260 746
rect 219 736 220 740
rect -4 722 -1 726
rect 408 740 409 744
rect 329 734 330 738
rect 105 719 106 723
rect -82 706 -81 710
rect -204 682 -203 686
rect -208 646 -203 682
rect -201 646 -197 686
rect -195 650 -190 686
rect -182 682 -181 686
rect -186 666 -181 682
rect -179 670 -174 686
rect -179 666 -178 670
rect -166 682 -165 686
rect -170 666 -165 682
rect -163 670 -158 686
rect -163 666 -162 670
rect -120 678 -119 682
rect -124 662 -119 678
rect -117 666 -110 682
rect 27 694 28 698
rect -117 662 -114 666
rect 23 658 28 694
rect 30 658 38 698
rect 40 662 45 698
rect 101 703 106 719
rect 108 707 113 723
rect 325 718 330 734
rect 332 722 337 738
rect 404 724 409 740
rect 411 728 416 744
rect 411 724 412 728
rect 332 718 333 722
rect 108 703 109 707
rect 470 685 471 689
rect 40 658 41 662
rect -195 646 -194 650
rect 96 657 97 661
rect 92 621 97 657
rect 99 621 107 661
rect 109 625 114 661
rect 438 656 439 660
rect 359 650 360 654
rect 319 644 320 648
rect 109 621 110 625
rect 131 637 132 641
rect 127 621 132 637
rect 134 625 139 641
rect 315 628 320 644
rect 322 632 327 648
rect 355 634 360 650
rect 362 638 367 654
rect 362 634 363 638
rect 398 650 399 654
rect 394 634 399 650
rect 401 638 406 654
rect 434 640 439 656
rect 441 644 446 660
rect 466 649 471 685
rect 473 649 477 689
rect 479 653 484 689
rect 492 685 493 689
rect 488 669 493 685
rect 495 673 500 689
rect 495 669 496 673
rect 508 685 509 689
rect 504 669 509 685
rect 511 673 516 689
rect 511 669 512 673
rect 554 681 555 685
rect 550 665 555 681
rect 557 669 564 685
rect 557 665 560 669
rect 479 649 480 653
rect 441 640 442 644
rect 401 634 402 638
rect 322 628 323 632
rect 134 621 135 625
rect -101 603 -100 607
rect -105 567 -100 603
rect -98 567 -94 607
rect -92 571 -87 607
rect -79 603 -78 607
rect -83 587 -78 603
rect -76 591 -71 607
rect -76 587 -75 591
rect -63 603 -62 607
rect -67 587 -62 603
rect -60 591 -55 607
rect -60 587 -59 591
rect -17 599 -16 603
rect -21 583 -16 599
rect -14 587 -7 603
rect 162 612 163 616
rect -14 583 -11 587
rect 158 596 163 612
rect 165 600 173 616
rect 165 596 167 600
rect 171 596 173 600
rect 175 612 176 616
rect 175 596 180 612
rect -92 567 -91 571
rect -212 541 -211 545
rect -216 505 -211 541
rect -209 505 -205 545
rect -203 509 -198 545
rect -190 541 -189 545
rect -194 525 -189 541
rect -187 529 -182 545
rect -187 525 -186 529
rect -174 541 -173 545
rect -178 525 -173 541
rect -171 529 -166 545
rect -171 525 -170 529
rect -128 537 -127 541
rect -132 521 -127 537
rect -125 525 -118 541
rect 23 562 28 578
rect 27 558 28 562
rect 30 574 32 578
rect 36 574 38 578
rect 30 558 38 574
rect 40 562 45 578
rect 40 558 41 562
rect 96 559 97 563
rect -125 521 -122 525
rect -203 505 -202 509
rect 22 520 23 524
rect 18 484 23 520
rect 25 484 33 524
rect 35 488 40 524
rect 92 523 97 559
rect 99 523 107 563
rect 109 527 114 563
rect 327 562 328 566
rect 323 546 328 562
rect 330 550 335 566
rect 330 546 331 550
rect 418 562 419 566
rect 414 546 419 562
rect 421 550 426 566
rect 421 546 422 550
rect 109 523 110 527
rect 154 527 155 531
rect 150 511 155 527
rect 157 515 165 531
rect 157 511 159 515
rect 163 511 165 515
rect 167 527 168 531
rect 167 511 172 527
rect 188 527 189 531
rect 184 511 189 527
rect 191 515 196 531
rect 191 511 192 515
rect 35 484 36 488
rect 86 469 87 473
rect -103 442 -102 446
rect -107 406 -102 442
rect -100 406 -96 446
rect -94 410 -89 446
rect -81 442 -80 446
rect -85 426 -80 442
rect -78 430 -73 446
rect -78 426 -77 430
rect -65 442 -64 446
rect -69 426 -64 442
rect -62 430 -57 446
rect -62 426 -61 430
rect -19 438 -18 442
rect -23 422 -18 438
rect -16 426 -9 442
rect -16 422 -13 426
rect 82 433 87 469
rect 89 433 97 473
rect 99 437 104 473
rect 482 507 483 511
rect 357 478 358 482
rect 317 472 318 476
rect 209 464 210 468
rect 99 433 100 437
rect 121 449 122 453
rect 117 433 122 449
rect 124 437 129 453
rect 124 433 125 437
rect -94 406 -93 410
rect -227 388 -226 392
rect -231 352 -226 388
rect -224 352 -220 392
rect -218 356 -213 392
rect -205 388 -204 392
rect -209 372 -204 388
rect -202 376 -197 392
rect -202 372 -201 376
rect -189 388 -188 392
rect -193 372 -188 388
rect -186 376 -181 392
rect -186 372 -185 376
rect -143 384 -142 388
rect -147 368 -142 384
rect -140 372 -133 388
rect -140 368 -137 372
rect 159 425 160 429
rect 155 409 160 425
rect 162 413 170 429
rect 162 409 164 413
rect 168 409 170 413
rect 172 425 173 429
rect 205 428 210 464
rect 212 428 220 468
rect 222 432 227 468
rect 313 456 318 472
rect 320 460 325 476
rect 353 462 358 478
rect 360 466 365 482
rect 448 478 449 482
rect 360 462 361 466
rect 408 472 409 476
rect 320 456 321 460
rect 222 428 223 432
rect 244 444 245 448
rect 240 428 245 444
rect 247 432 252 448
rect 404 456 409 472
rect 411 460 416 476
rect 444 462 449 478
rect 451 466 456 482
rect 478 471 483 507
rect 485 471 489 511
rect 491 475 496 511
rect 504 507 505 511
rect 500 491 505 507
rect 507 495 512 511
rect 507 491 508 495
rect 520 507 521 511
rect 516 491 521 507
rect 523 495 528 511
rect 523 491 524 495
rect 566 503 567 507
rect 562 487 567 503
rect 569 491 576 507
rect 569 487 572 491
rect 491 471 492 475
rect 451 462 452 466
rect 411 456 412 460
rect 247 428 248 432
rect 172 409 177 425
rect 18 388 23 404
rect 22 384 23 388
rect 25 400 27 404
rect 31 400 33 404
rect 25 384 33 400
rect 35 388 40 404
rect 332 396 333 400
rect 35 384 36 388
rect 77 371 78 375
rect -218 352 -217 356
rect 21 347 22 351
rect 17 311 22 347
rect 24 311 32 351
rect 34 315 39 351
rect 73 335 78 371
rect 80 335 88 375
rect 90 339 95 375
rect 328 380 333 396
rect 335 384 340 400
rect 335 380 336 384
rect 419 396 420 400
rect 415 380 420 396
rect 422 384 427 400
rect 422 380 423 384
rect 90 335 91 339
rect 198 332 199 336
rect 34 311 35 315
rect 194 316 199 332
rect 201 320 209 336
rect 201 316 203 320
rect 207 316 209 320
rect 211 332 212 336
rect 211 316 216 332
rect 232 332 233 336
rect 228 316 233 332
rect 235 320 240 336
rect 482 350 483 354
rect 235 316 236 320
rect 362 312 363 316
rect 322 306 323 310
rect 84 278 85 282
rect -110 269 -109 273
rect -114 233 -109 269
rect -107 233 -103 273
rect -101 237 -96 273
rect -88 269 -87 273
rect -92 253 -87 269
rect -85 257 -80 273
rect -85 253 -84 257
rect -72 269 -71 273
rect -76 253 -71 269
rect -69 257 -64 273
rect -69 253 -68 257
rect -26 265 -25 269
rect -30 249 -25 265
rect -23 253 -16 269
rect -23 249 -20 253
rect -101 233 -100 237
rect 80 242 85 278
rect 87 242 95 282
rect 97 246 102 282
rect 318 290 323 306
rect 325 294 330 310
rect 358 296 363 312
rect 365 300 370 316
rect 449 312 450 316
rect 365 296 366 300
rect 409 306 410 310
rect 325 290 326 294
rect 405 290 410 306
rect 412 294 417 310
rect 445 296 450 312
rect 452 300 457 316
rect 478 314 483 350
rect 485 314 489 354
rect 491 318 496 354
rect 504 350 505 354
rect 500 334 505 350
rect 507 338 512 354
rect 507 334 508 338
rect 520 350 521 354
rect 516 334 521 350
rect 523 338 528 354
rect 523 334 524 338
rect 566 346 567 350
rect 562 330 567 346
rect 569 334 576 350
rect 569 330 572 334
rect 491 314 492 318
rect 452 296 453 300
rect 412 290 413 294
rect 97 242 98 246
rect 119 258 120 262
rect 115 242 120 258
rect 122 246 127 262
rect 122 242 123 246
rect 204 247 205 251
rect 17 215 22 231
rect 21 211 22 215
rect 24 227 26 231
rect 30 227 32 231
rect 24 211 32 227
rect 34 215 39 231
rect 159 233 160 237
rect 34 211 35 215
rect 155 217 160 233
rect 162 221 170 237
rect 162 217 164 221
rect 168 217 170 221
rect 172 233 173 237
rect 172 217 177 233
rect 200 211 205 247
rect 207 211 215 251
rect 217 215 222 251
rect 416 233 417 237
rect 217 211 218 215
rect 239 227 240 231
rect 235 211 240 227
rect 242 215 247 231
rect 412 217 417 233
rect 419 221 424 237
rect 419 217 420 221
rect 482 231 483 235
rect 242 211 243 215
rect 84 180 85 184
rect -228 158 -227 162
rect -232 122 -227 158
rect -225 122 -221 162
rect -219 126 -214 162
rect -206 158 -205 162
rect -210 142 -205 158
rect -203 146 -198 162
rect -203 142 -202 146
rect -190 158 -189 162
rect -194 142 -189 158
rect -187 146 -182 162
rect -187 142 -186 146
rect -144 154 -143 158
rect -148 138 -143 154
rect -141 142 -134 158
rect -141 138 -138 142
rect 23 147 24 151
rect -219 122 -218 126
rect 19 111 24 147
rect 26 111 34 151
rect 36 115 41 151
rect 80 144 85 180
rect 87 144 95 184
rect 97 148 102 184
rect 478 195 483 231
rect 485 195 489 235
rect 491 199 496 235
rect 504 231 505 235
rect 500 215 505 231
rect 507 219 512 235
rect 507 215 508 219
rect 520 231 521 235
rect 516 215 521 231
rect 523 219 528 235
rect 523 215 524 219
rect 566 227 567 231
rect 562 211 567 227
rect 569 215 576 231
rect 569 211 572 215
rect 491 195 492 199
rect 334 191 335 195
rect 330 175 335 191
rect 337 179 342 195
rect 337 175 338 179
rect 97 144 98 148
rect 161 148 162 152
rect 157 132 162 148
rect 164 136 172 152
rect 164 132 166 136
rect 170 132 172 136
rect 174 148 175 152
rect 174 132 179 148
rect 195 148 196 152
rect 191 132 196 148
rect 198 136 203 152
rect 446 149 447 153
rect 198 132 199 136
rect 36 111 37 115
rect 406 143 407 147
rect 402 127 407 143
rect 409 131 414 147
rect 442 133 447 149
rect 449 137 454 153
rect 449 133 450 137
rect 409 127 410 131
rect 78 90 79 94
rect -113 71 -112 75
rect -117 35 -112 71
rect -110 35 -106 75
rect -104 39 -99 75
rect -91 71 -90 75
rect -95 55 -90 71
rect -88 59 -83 75
rect -88 55 -87 59
rect -75 71 -74 75
rect -79 55 -74 71
rect -72 59 -67 75
rect -72 55 -71 59
rect -29 67 -28 71
rect -33 51 -28 67
rect -26 55 -19 71
rect -26 51 -23 55
rect 74 54 79 90
rect 81 54 89 94
rect 91 58 96 94
rect 364 107 365 111
rect 324 101 325 105
rect 220 95 221 99
rect 91 54 92 58
rect 113 70 114 74
rect 109 54 114 70
rect 116 58 121 74
rect 116 54 117 58
rect 137 69 138 73
rect -104 35 -103 39
rect 133 53 138 69
rect 140 57 148 73
rect 140 53 142 57
rect 146 53 148 57
rect 150 69 151 73
rect 150 53 155 69
rect 216 59 221 95
rect 223 59 231 99
rect 233 63 238 99
rect 320 85 325 101
rect 327 89 332 105
rect 360 91 365 107
rect 367 95 372 111
rect 485 108 486 112
rect 367 91 368 95
rect 327 85 328 89
rect 233 59 234 63
rect 255 75 256 79
rect 251 59 256 75
rect 258 63 263 79
rect 258 59 259 63
rect 481 72 486 108
rect 488 72 492 112
rect 494 76 499 112
rect 507 108 508 112
rect 503 92 508 108
rect 510 96 515 112
rect 510 92 511 96
rect 523 108 524 112
rect 519 92 524 108
rect 526 96 531 112
rect 526 92 527 96
rect 569 104 570 108
rect 565 88 570 104
rect 572 92 579 108
rect 572 88 575 92
rect 494 72 495 76
rect 19 15 24 31
rect 23 11 24 15
rect 26 27 28 31
rect 32 27 34 31
rect 26 11 34 27
rect 36 15 41 31
rect 36 11 37 15
<< ndcontact >>
rect -63 817 -59 821
rect -95 795 -91 799
rect -87 801 -83 805
rect -41 817 -37 821
rect -11 809 -7 813
rect -1 815 3 819
rect -19 801 -15 805
rect 222 804 226 808
rect 230 810 234 814
rect 340 804 344 808
rect -49 781 -45 785
rect 216 772 220 776
rect 308 782 312 786
rect 316 788 320 792
rect 245 775 249 779
rect 362 804 366 808
rect 392 796 396 800
rect 402 802 406 806
rect 384 788 388 792
rect 354 768 358 772
rect -63 706 -59 710
rect -95 684 -91 688
rect -87 690 -83 694
rect -41 706 -37 710
rect -11 698 -7 702
rect -1 704 3 708
rect -19 690 -15 694
rect -49 670 -45 674
rect 60 696 64 700
rect 78 712 82 716
rect 212 714 216 718
rect 220 720 224 724
rect 252 710 256 714
rect 260 726 264 730
rect 325 696 329 700
rect 333 702 337 706
rect 404 702 408 706
rect 412 708 416 712
rect 101 681 105 685
rect 109 687 113 691
rect 319 664 323 668
rect 348 667 352 671
rect 398 670 402 674
rect 427 673 431 677
rect -176 646 -172 650
rect -208 624 -204 628
rect -200 630 -196 634
rect -154 646 -150 650
rect -124 638 -120 642
rect -114 644 -110 648
rect -132 630 -128 634
rect 23 629 27 633
rect 32 635 36 639
rect 41 629 45 633
rect 498 649 502 653
rect -162 610 -158 614
rect 23 614 27 618
rect 41 598 45 602
rect 92 593 96 597
rect 101 599 105 603
rect 127 597 131 601
rect 135 603 139 607
rect 110 593 114 597
rect 315 606 319 610
rect 323 612 327 616
rect 355 602 359 606
rect 363 618 367 622
rect 394 612 398 616
rect 402 618 406 622
rect 434 608 438 612
rect 442 624 446 628
rect 466 627 470 631
rect 474 633 478 637
rect 520 649 524 653
rect 550 641 554 645
rect 560 647 564 651
rect 542 633 546 637
rect 512 613 516 617
rect -73 567 -69 571
rect -105 545 -101 549
rect -97 551 -93 555
rect -51 567 -47 571
rect -21 559 -17 563
rect -11 565 -7 569
rect -29 551 -25 555
rect -59 531 -55 535
rect -184 505 -180 509
rect -216 483 -212 487
rect -208 489 -204 493
rect -162 505 -158 509
rect -132 497 -128 501
rect -122 503 -118 507
rect -140 489 -136 493
rect 158 557 162 561
rect 176 573 180 577
rect 323 524 327 528
rect 331 530 335 534
rect 414 524 418 528
rect 422 530 426 534
rect 92 495 96 499
rect 101 501 105 505
rect 110 495 114 499
rect -170 469 -166 473
rect 18 455 22 459
rect 27 461 31 465
rect 36 455 40 459
rect 18 440 22 444
rect 150 472 154 476
rect 168 488 172 492
rect 184 489 188 493
rect 192 495 196 499
rect 317 492 321 496
rect 346 495 350 499
rect 408 492 412 496
rect 437 495 441 499
rect 36 424 40 428
rect -75 406 -71 410
rect -107 384 -103 388
rect -99 390 -95 394
rect -53 406 -49 410
rect -23 398 -19 402
rect -13 404 -9 408
rect 82 405 86 409
rect 91 411 95 415
rect 117 409 121 413
rect 125 415 129 419
rect 510 471 514 475
rect 313 434 317 438
rect 321 440 325 444
rect 353 430 357 434
rect 361 446 365 450
rect 404 434 408 438
rect 412 440 416 444
rect 444 430 448 434
rect 452 446 456 450
rect 478 449 482 453
rect 486 455 490 459
rect 532 471 536 475
rect 562 463 566 467
rect 572 469 576 473
rect 554 455 558 459
rect 524 435 528 439
rect 100 405 104 409
rect -31 390 -27 394
rect 205 400 209 404
rect 214 406 218 410
rect 240 404 244 408
rect 248 410 252 414
rect 223 400 227 404
rect -61 370 -57 374
rect -199 352 -195 356
rect -231 330 -227 334
rect -223 336 -219 340
rect -177 352 -173 356
rect -147 344 -143 348
rect -137 350 -133 354
rect -155 336 -151 340
rect -185 316 -181 320
rect 155 370 159 374
rect 173 386 177 390
rect 328 358 332 362
rect 336 364 340 368
rect 415 358 419 362
rect 423 364 427 368
rect 73 307 77 311
rect 82 313 86 317
rect 322 326 326 330
rect 351 329 355 333
rect 409 326 413 330
rect 438 329 442 333
rect 91 307 95 311
rect 17 282 21 286
rect 26 288 30 292
rect 35 282 39 286
rect 17 267 21 271
rect 35 251 39 255
rect -82 233 -78 237
rect -114 211 -110 215
rect -106 217 -102 221
rect -60 233 -56 237
rect -30 225 -26 229
rect -20 231 -16 235
rect 194 277 198 281
rect 212 293 216 297
rect 228 294 232 298
rect 236 300 240 304
rect 510 314 514 318
rect 318 268 322 272
rect 326 274 330 278
rect 358 264 362 268
rect 366 280 370 284
rect 478 292 482 296
rect 486 298 490 302
rect 405 268 409 272
rect 413 274 417 278
rect 445 264 449 268
rect 453 280 457 284
rect 532 314 536 318
rect 562 306 566 310
rect 572 312 576 316
rect 554 298 558 302
rect 524 278 528 282
rect -38 217 -34 221
rect 80 214 84 218
rect 89 220 93 224
rect 115 218 119 222
rect 123 224 127 228
rect 98 214 102 218
rect -68 197 -64 201
rect -200 122 -196 126
rect -232 100 -228 104
rect -224 106 -220 110
rect -178 122 -174 126
rect -148 114 -144 118
rect -138 120 -134 124
rect 155 178 159 182
rect 173 194 177 198
rect 200 183 204 187
rect 209 189 213 193
rect 235 187 239 191
rect 243 193 247 197
rect 412 195 416 199
rect 420 201 424 205
rect 510 195 514 199
rect 218 183 222 187
rect 406 163 410 167
rect 478 173 482 177
rect 486 179 490 183
rect 435 166 439 170
rect 330 153 334 157
rect 338 159 342 163
rect 532 195 536 199
rect 562 187 566 191
rect 572 193 576 197
rect 554 179 558 183
rect 524 159 528 163
rect 80 116 84 120
rect 89 122 93 126
rect 98 116 102 120
rect 324 121 328 125
rect 353 124 357 128
rect -156 106 -152 110
rect -186 86 -182 90
rect 19 82 23 86
rect 28 88 32 92
rect 37 82 41 86
rect 19 67 23 71
rect 37 51 41 55
rect 157 93 161 97
rect 175 109 179 113
rect 191 110 195 114
rect 199 116 203 120
rect -85 35 -81 39
rect -117 13 -113 17
rect -109 19 -105 23
rect -63 35 -59 39
rect -33 27 -29 31
rect -23 33 -19 37
rect 402 105 406 109
rect 410 111 414 115
rect 442 101 446 105
rect 450 117 454 121
rect 320 63 324 67
rect 328 69 332 73
rect 360 59 364 63
rect 368 75 372 79
rect 513 72 517 76
rect -41 19 -37 23
rect 74 26 78 30
rect 83 32 87 36
rect 109 30 113 34
rect 117 36 121 40
rect 481 50 485 54
rect 489 56 493 60
rect 92 26 96 30
rect 133 14 137 18
rect 151 30 155 34
rect 216 31 220 35
rect 225 37 229 41
rect 251 35 255 39
rect 259 41 263 45
rect 535 72 539 76
rect 565 64 569 68
rect 575 70 579 74
rect 557 56 561 60
rect 527 36 531 40
rect 234 31 238 35
rect -71 -1 -67 3
<< pdcontact >>
rect -95 853 -91 857
rect -73 853 -69 857
rect -65 837 -61 841
rect -57 853 -53 857
rect -49 837 -45 841
rect -11 849 -7 853
rect -1 833 3 837
rect 222 842 226 846
rect 230 826 234 830
rect 308 840 312 844
rect -81 817 -77 821
rect 330 840 334 844
rect 338 824 342 828
rect 346 840 350 844
rect 354 824 358 828
rect 392 836 396 840
rect 402 820 406 824
rect 322 804 326 808
rect 252 758 256 762
rect 60 751 64 755
rect -95 742 -91 746
rect -73 742 -69 746
rect -65 726 -61 730
rect -57 742 -53 746
rect -49 726 -45 730
rect -11 738 -7 742
rect 69 735 73 739
rect 78 751 82 755
rect 212 752 216 756
rect 260 742 264 746
rect 220 736 224 740
rect -1 722 3 726
rect 404 740 408 744
rect 325 734 329 738
rect 101 719 105 723
rect -81 706 -77 710
rect -208 682 -204 686
rect -186 682 -182 686
rect -178 666 -174 670
rect -170 682 -166 686
rect -162 666 -158 670
rect -124 678 -120 682
rect 23 694 27 698
rect -114 662 -110 666
rect 412 724 416 728
rect 333 718 337 722
rect 109 703 113 707
rect 466 685 470 689
rect 41 658 45 662
rect -194 646 -190 650
rect 92 657 96 661
rect 434 656 438 660
rect 355 650 359 654
rect 315 644 319 648
rect 110 621 114 625
rect 127 637 131 641
rect 363 634 367 638
rect 394 650 398 654
rect 488 685 492 689
rect 496 669 500 673
rect 504 685 508 689
rect 512 669 516 673
rect 550 681 554 685
rect 560 665 564 669
rect 480 649 484 653
rect 442 640 446 644
rect 402 634 406 638
rect 323 628 327 632
rect 135 621 139 625
rect -105 603 -101 607
rect -83 603 -79 607
rect -75 587 -71 591
rect -67 603 -63 607
rect -59 587 -55 591
rect -21 599 -17 603
rect 158 612 162 616
rect -11 583 -7 587
rect 167 596 171 600
rect 176 612 180 616
rect -91 567 -87 571
rect -216 541 -212 545
rect -194 541 -190 545
rect -186 525 -182 529
rect -178 541 -174 545
rect -170 525 -166 529
rect -132 537 -128 541
rect 23 558 27 562
rect 32 574 36 578
rect 41 558 45 562
rect 92 559 96 563
rect -122 521 -118 525
rect -202 505 -198 509
rect 18 520 22 524
rect 323 562 327 566
rect 331 546 335 550
rect 414 562 418 566
rect 422 546 426 550
rect 110 523 114 527
rect 150 527 154 531
rect 159 511 163 515
rect 168 527 172 531
rect 184 527 188 531
rect 192 511 196 515
rect 36 484 40 488
rect 82 469 86 473
rect -107 442 -103 446
rect -85 442 -81 446
rect -77 426 -73 430
rect -69 442 -65 446
rect -61 426 -57 430
rect -23 438 -19 442
rect -13 422 -9 426
rect 478 507 482 511
rect 353 478 357 482
rect 313 472 317 476
rect 205 464 209 468
rect 100 433 104 437
rect 117 449 121 453
rect 125 433 129 437
rect -93 406 -89 410
rect -231 388 -227 392
rect -209 388 -205 392
rect -201 372 -197 376
rect -193 388 -189 392
rect -185 372 -181 376
rect -147 384 -143 388
rect -137 368 -133 372
rect 155 425 159 429
rect 164 409 168 413
rect 173 425 177 429
rect 444 478 448 482
rect 361 462 365 466
rect 404 472 408 476
rect 321 456 325 460
rect 223 428 227 432
rect 240 444 244 448
rect 500 507 504 511
rect 508 491 512 495
rect 516 507 520 511
rect 524 491 528 495
rect 562 503 566 507
rect 572 487 576 491
rect 492 471 496 475
rect 452 462 456 466
rect 412 456 416 460
rect 248 428 252 432
rect 18 384 22 388
rect 27 400 31 404
rect 328 396 332 400
rect 36 384 40 388
rect 73 371 77 375
rect -217 352 -213 356
rect 17 347 21 351
rect 336 380 340 384
rect 415 396 419 400
rect 423 380 427 384
rect 91 335 95 339
rect 194 332 198 336
rect 35 311 39 315
rect 203 316 207 320
rect 212 332 216 336
rect 228 332 232 336
rect 478 350 482 354
rect 236 316 240 320
rect 358 312 362 316
rect 318 306 322 310
rect 80 278 84 282
rect -114 269 -110 273
rect -92 269 -88 273
rect -84 253 -80 257
rect -76 269 -72 273
rect -68 253 -64 257
rect -30 265 -26 269
rect -20 249 -16 253
rect -100 233 -96 237
rect 445 312 449 316
rect 366 296 370 300
rect 405 306 409 310
rect 326 290 330 294
rect 500 350 504 354
rect 508 334 512 338
rect 516 350 520 354
rect 524 334 528 338
rect 562 346 566 350
rect 572 330 576 334
rect 492 314 496 318
rect 453 296 457 300
rect 413 290 417 294
rect 98 242 102 246
rect 115 258 119 262
rect 123 242 127 246
rect 200 247 204 251
rect 17 211 21 215
rect 26 227 30 231
rect 155 233 159 237
rect 35 211 39 215
rect 164 217 168 221
rect 173 233 177 237
rect 412 233 416 237
rect 218 211 222 215
rect 235 227 239 231
rect 420 217 424 221
rect 478 231 482 235
rect 243 211 247 215
rect 80 180 84 184
rect -232 158 -228 162
rect -210 158 -206 162
rect -202 142 -198 146
rect -194 158 -190 162
rect -186 142 -182 146
rect -148 154 -144 158
rect -138 138 -134 142
rect 19 147 23 151
rect -218 122 -214 126
rect 500 231 504 235
rect 508 215 512 219
rect 516 231 520 235
rect 524 215 528 219
rect 562 227 566 231
rect 572 211 576 215
rect 492 195 496 199
rect 330 191 334 195
rect 338 175 342 179
rect 98 144 102 148
rect 157 148 161 152
rect 166 132 170 136
rect 175 148 179 152
rect 191 148 195 152
rect 442 149 446 153
rect 199 132 203 136
rect 37 111 41 115
rect 402 143 406 147
rect 450 133 454 137
rect 410 127 414 131
rect 74 90 78 94
rect -117 71 -113 75
rect -95 71 -91 75
rect -87 55 -83 59
rect -79 71 -75 75
rect -71 55 -67 59
rect -33 67 -29 71
rect -23 51 -19 55
rect 360 107 364 111
rect 320 101 324 105
rect 216 95 220 99
rect 92 54 96 58
rect 109 70 113 74
rect 117 54 121 58
rect 133 69 137 73
rect -103 35 -99 39
rect 142 53 146 57
rect 151 69 155 73
rect 481 108 485 112
rect 368 91 372 95
rect 328 85 332 89
rect 234 59 238 63
rect 251 75 255 79
rect 259 59 263 63
rect 503 108 507 112
rect 511 92 515 96
rect 519 108 523 112
rect 527 92 531 96
rect 565 104 569 108
rect 575 88 579 92
rect 495 72 499 76
rect 19 11 23 15
rect 28 27 32 31
rect 37 11 41 15
<< polysilicon >>
rect -90 857 -88 860
rect -84 857 -82 864
rect -68 857 -66 869
rect -52 857 -50 860
rect -6 853 -4 861
rect -68 834 -66 837
rect -52 832 -50 837
rect 227 846 229 849
rect -58 821 -56 824
rect -6 826 -4 833
rect 313 844 315 847
rect 319 844 321 851
rect 335 844 337 856
rect 351 844 353 847
rect -52 821 -50 822
rect -34 821 -32 822
rect -25 821 -23 824
rect -90 805 -88 817
rect -84 814 -82 817
rect -90 792 -88 795
rect -6 819 -4 822
rect 227 814 229 826
rect -6 806 -4 809
rect 397 840 399 848
rect 335 821 337 824
rect 351 819 353 824
rect 345 808 347 811
rect 397 813 399 820
rect 351 808 353 809
rect 369 808 371 809
rect 378 808 380 811
rect 227 801 229 804
rect -34 798 -32 801
rect -25 798 -23 801
rect 242 795 244 796
rect 213 792 215 793
rect -58 780 -56 781
rect -52 778 -50 781
rect 313 792 315 804
rect 319 801 321 804
rect 313 779 315 782
rect 242 772 244 775
rect 213 769 215 772
rect 397 806 399 809
rect 397 793 399 796
rect 369 785 371 788
rect 378 785 380 788
rect 345 767 347 768
rect 257 762 259 765
rect 351 765 353 768
rect -90 746 -88 749
rect -84 746 -82 753
rect -68 746 -66 758
rect 65 755 67 759
rect 75 755 77 759
rect 217 756 219 759
rect -52 746 -50 749
rect -6 742 -4 750
rect -68 723 -66 726
rect -52 721 -50 726
rect 409 744 411 747
rect -58 710 -56 713
rect -6 715 -4 722
rect 65 716 67 735
rect 75 716 77 735
rect 106 723 108 726
rect 217 724 219 736
rect 257 730 259 742
rect 330 738 332 741
rect -52 710 -50 711
rect -34 710 -32 711
rect -25 710 -23 713
rect -203 686 -201 689
rect -197 686 -195 693
rect -181 686 -179 698
rect -90 694 -88 706
rect -84 703 -82 706
rect -165 686 -163 689
rect -119 682 -117 690
rect -181 663 -179 666
rect -165 661 -163 666
rect -90 681 -88 684
rect -6 708 -4 711
rect 28 698 30 701
rect 38 698 40 701
rect -6 695 -4 698
rect -34 687 -32 690
rect -25 687 -23 690
rect -58 669 -56 670
rect -52 667 -50 670
rect -171 650 -169 653
rect -119 655 -117 662
rect 217 711 219 714
rect 257 707 259 710
rect 330 706 332 718
rect 409 712 411 724
rect 65 693 67 696
rect 75 693 77 696
rect 106 691 108 703
rect 409 699 411 702
rect 330 693 332 696
rect 424 693 426 694
rect 395 690 397 691
rect 345 687 347 688
rect 316 684 318 685
rect 106 678 108 681
rect 471 689 473 692
rect 477 689 479 696
rect 493 689 495 701
rect 509 689 511 692
rect 424 670 426 673
rect 395 667 397 670
rect 345 664 347 667
rect 97 661 99 664
rect 107 661 109 664
rect 316 661 318 664
rect -165 650 -163 651
rect -147 650 -145 651
rect -138 650 -136 653
rect -203 634 -201 646
rect -197 643 -195 646
rect -203 621 -201 624
rect -119 648 -117 651
rect 28 639 30 658
rect 38 639 40 658
rect -119 635 -117 638
rect -147 627 -145 630
rect -138 627 -136 630
rect 28 626 30 629
rect 38 626 40 629
rect 439 660 441 663
rect 360 654 362 657
rect 399 654 401 657
rect 320 648 322 651
rect 132 641 134 644
rect 555 685 557 693
rect 493 666 495 669
rect 509 664 511 669
rect 503 653 505 656
rect 555 658 557 665
rect 509 653 511 654
rect 527 653 529 654
rect 536 653 538 656
rect -171 609 -169 610
rect -165 607 -163 610
rect -100 607 -98 610
rect -94 607 -92 614
rect -78 607 -76 619
rect 28 618 30 621
rect 38 618 40 621
rect -62 607 -60 610
rect -16 603 -14 611
rect -78 584 -76 587
rect -62 582 -60 587
rect 97 603 99 621
rect 107 603 109 621
rect 132 607 134 621
rect 163 616 165 620
rect 173 616 175 620
rect 320 616 322 628
rect 360 622 362 634
rect 399 622 401 634
rect 439 628 441 640
rect 471 637 473 649
rect 477 646 479 649
rect -68 571 -66 574
rect -16 576 -14 583
rect 28 578 30 598
rect 38 578 40 598
rect 132 594 134 597
rect 320 603 322 606
rect 399 609 401 612
rect 471 624 473 627
rect 555 651 557 654
rect 555 638 557 641
rect 527 630 529 633
rect 536 630 538 633
rect 503 612 505 613
rect 509 610 511 613
rect 439 605 441 608
rect 360 599 362 602
rect 97 590 99 593
rect 107 590 109 593
rect -62 571 -60 572
rect -44 571 -42 572
rect -35 571 -33 574
rect -211 545 -209 548
rect -205 545 -203 552
rect -189 545 -187 557
rect -100 555 -98 567
rect -94 564 -92 567
rect -173 545 -171 548
rect -127 541 -125 549
rect -100 542 -98 545
rect -189 522 -187 525
rect -173 520 -171 525
rect -16 569 -14 572
rect -16 556 -14 559
rect 163 577 165 596
rect 173 577 175 596
rect 97 563 99 566
rect 107 563 109 566
rect 28 554 30 558
rect 38 554 40 558
rect -44 548 -42 551
rect -35 548 -33 551
rect -68 530 -66 531
rect -62 528 -60 531
rect 23 524 25 527
rect 33 524 35 527
rect -179 509 -177 512
rect -127 514 -125 521
rect -173 509 -171 510
rect -155 509 -153 510
rect -146 509 -144 512
rect -211 493 -209 505
rect -205 502 -203 505
rect -211 480 -209 483
rect -127 507 -125 510
rect -127 494 -125 497
rect -155 486 -153 489
rect -146 486 -144 489
rect 328 566 330 569
rect 419 566 421 569
rect 163 554 165 557
rect 173 554 175 557
rect 155 531 157 535
rect 165 531 167 535
rect 328 534 330 546
rect 419 534 421 546
rect 189 531 191 534
rect 97 505 99 523
rect 107 505 109 523
rect 328 521 330 524
rect 419 521 421 524
rect 343 515 345 516
rect 314 512 316 513
rect 97 492 99 495
rect 107 492 109 495
rect 155 492 157 511
rect 165 492 167 511
rect 189 499 191 511
rect -179 468 -177 469
rect -173 466 -171 469
rect 23 465 25 484
rect 33 465 35 484
rect 87 473 89 476
rect 97 473 99 476
rect -102 446 -100 449
rect -96 446 -94 453
rect -80 446 -78 458
rect 23 452 25 455
rect 33 452 35 455
rect -64 446 -62 449
rect -18 442 -16 450
rect 23 444 25 447
rect 33 444 35 447
rect -80 423 -78 426
rect -64 421 -62 426
rect 434 515 436 516
rect 405 512 407 513
rect 343 492 345 495
rect 483 511 485 514
rect 489 511 491 518
rect 505 511 507 523
rect 521 511 523 514
rect 434 492 436 495
rect 314 489 316 492
rect 405 489 407 492
rect 189 486 191 489
rect 358 482 360 485
rect 449 482 451 485
rect 318 476 320 479
rect 155 469 157 472
rect 165 469 167 472
rect 210 468 212 471
rect 220 468 222 471
rect 122 453 124 456
rect -70 410 -68 413
rect -18 415 -16 422
rect -64 410 -62 411
rect -46 410 -44 411
rect -37 410 -35 413
rect -226 392 -224 395
rect -220 392 -218 399
rect -204 392 -202 404
rect -188 392 -186 395
rect -142 388 -140 396
rect -102 394 -100 406
rect -96 403 -94 406
rect -204 369 -202 372
rect -188 367 -186 372
rect -102 381 -100 384
rect -18 408 -16 411
rect 23 404 25 424
rect 33 404 35 424
rect 87 415 89 433
rect 97 415 99 433
rect 122 419 124 433
rect 160 429 162 433
rect 170 429 172 433
rect 409 476 411 479
rect 245 448 247 451
rect 318 444 320 456
rect 358 450 360 462
rect 567 507 569 515
rect 505 488 507 491
rect 521 486 523 491
rect 515 475 517 478
rect 567 480 569 487
rect 521 475 523 476
rect 539 475 541 476
rect 548 475 550 478
rect 318 431 320 434
rect 409 444 411 456
rect 449 450 451 462
rect 483 459 485 471
rect 489 468 491 471
rect 409 431 411 434
rect 483 446 485 449
rect 567 473 569 476
rect 567 460 569 463
rect 539 452 541 455
rect 548 452 550 455
rect 515 434 517 435
rect 521 432 523 435
rect 210 410 212 428
rect 220 410 222 428
rect 245 414 247 428
rect 358 427 360 430
rect 449 427 451 430
rect 122 406 124 409
rect -18 395 -16 398
rect -46 387 -44 390
rect -37 387 -35 390
rect 87 402 89 405
rect 97 402 99 405
rect 160 390 162 409
rect 170 390 172 409
rect 245 401 247 404
rect 333 400 335 403
rect 420 400 422 403
rect 210 397 212 400
rect 220 397 222 400
rect 23 380 25 384
rect 33 380 35 384
rect 78 375 80 378
rect 88 375 90 378
rect -70 369 -68 370
rect -194 356 -192 359
rect -142 361 -140 368
rect -64 367 -62 370
rect -188 356 -186 357
rect -170 356 -168 357
rect -161 356 -159 359
rect -226 340 -224 352
rect -220 349 -218 352
rect -226 327 -224 330
rect -142 354 -140 357
rect 22 351 24 354
rect 32 351 34 354
rect -142 341 -140 344
rect -170 333 -168 336
rect -161 333 -159 336
rect -194 315 -192 316
rect -188 313 -186 316
rect 160 367 162 370
rect 170 367 172 370
rect 333 368 335 380
rect 420 368 422 380
rect 333 355 335 358
rect 420 355 422 358
rect 483 354 485 357
rect 489 354 491 361
rect 505 354 507 366
rect 521 354 523 357
rect 348 349 350 350
rect 319 346 321 347
rect 199 336 201 340
rect 209 336 211 340
rect 233 336 235 339
rect 78 317 80 335
rect 88 317 90 335
rect 22 292 24 311
rect 32 292 34 311
rect 435 349 437 350
rect 406 346 408 347
rect 348 326 350 329
rect 435 326 437 329
rect 319 323 321 326
rect 406 323 408 326
rect 363 316 365 319
rect 450 316 452 319
rect 78 304 80 307
rect 88 304 90 307
rect 199 297 201 316
rect 209 297 211 316
rect 233 304 235 316
rect 323 310 325 313
rect -109 273 -107 276
rect -103 273 -101 280
rect -87 273 -85 285
rect 85 282 87 285
rect 95 282 97 285
rect 22 279 24 282
rect 32 279 34 282
rect -71 273 -69 276
rect -25 269 -23 277
rect 22 271 24 274
rect 32 271 34 274
rect -87 250 -85 253
rect -71 248 -69 253
rect -77 237 -75 240
rect -25 242 -23 249
rect -71 237 -69 238
rect -53 237 -51 238
rect -44 237 -42 240
rect -109 221 -107 233
rect -103 230 -101 233
rect -109 208 -107 211
rect -25 235 -23 238
rect 22 231 24 251
rect 32 231 34 251
rect 233 291 235 294
rect 410 310 412 313
rect 323 278 325 290
rect 363 284 365 296
rect 567 350 569 358
rect 505 331 507 334
rect 521 329 523 334
rect 515 318 517 321
rect 567 323 569 330
rect 521 318 523 319
rect 539 318 541 319
rect 548 318 550 321
rect 483 302 485 314
rect 489 311 491 314
rect 199 274 201 277
rect 209 274 211 277
rect 323 265 325 268
rect 120 262 122 265
rect 410 278 412 290
rect 450 284 452 296
rect 483 289 485 292
rect 410 265 412 268
rect 567 316 569 319
rect 567 303 569 306
rect 539 295 541 298
rect 548 295 550 298
rect 515 277 517 278
rect 521 275 523 278
rect 363 261 365 264
rect 450 261 452 264
rect 205 251 207 254
rect 215 251 217 254
rect -25 222 -23 225
rect -53 214 -51 217
rect -44 214 -42 217
rect 85 224 87 242
rect 95 224 97 242
rect 120 228 122 242
rect 160 237 162 241
rect 170 237 172 241
rect 120 215 122 218
rect 85 211 87 214
rect 95 211 97 214
rect 22 207 24 211
rect 32 207 34 211
rect 160 198 162 217
rect 170 198 172 217
rect 417 237 419 240
rect 240 231 242 234
rect 483 235 485 238
rect 489 235 491 242
rect 505 235 507 247
rect 521 235 523 238
rect -77 196 -75 197
rect -71 194 -69 197
rect 85 184 87 187
rect 95 184 97 187
rect -227 162 -225 165
rect -221 162 -219 169
rect -205 162 -203 174
rect -189 162 -187 165
rect -143 158 -141 166
rect -205 139 -203 142
rect -189 137 -187 142
rect 24 151 26 154
rect 34 151 36 154
rect -195 126 -193 129
rect -143 131 -141 138
rect -189 126 -187 127
rect -171 126 -169 127
rect -162 126 -160 129
rect -227 110 -225 122
rect -221 119 -219 122
rect -227 97 -225 100
rect -143 124 -141 127
rect -143 111 -141 114
rect 205 193 207 211
rect 215 193 217 211
rect 240 197 242 211
rect 417 205 419 217
rect 335 195 337 198
rect 567 231 569 239
rect 505 212 507 215
rect 521 210 523 215
rect 515 199 517 202
rect 567 204 569 211
rect 521 199 523 200
rect 539 199 541 200
rect 548 199 550 202
rect 240 184 242 187
rect 205 180 207 183
rect 215 180 217 183
rect 160 175 162 178
rect 170 175 172 178
rect 417 192 419 195
rect 432 186 434 187
rect 403 183 405 184
rect 335 163 337 175
rect 483 183 485 195
rect 489 192 491 195
rect 483 170 485 173
rect 432 163 434 166
rect 162 152 164 156
rect 172 152 174 156
rect 196 152 198 155
rect 403 160 405 163
rect 567 197 569 200
rect 567 184 569 187
rect 539 176 541 179
rect 548 176 550 179
rect 515 158 517 159
rect 447 153 449 156
rect 521 156 523 159
rect 85 126 87 144
rect 95 126 97 144
rect 335 150 337 153
rect 407 147 409 150
rect 350 144 352 145
rect 321 141 323 142
rect 85 113 87 116
rect 95 113 97 116
rect 162 113 164 132
rect 172 113 174 132
rect 196 120 198 132
rect 350 121 352 124
rect -171 103 -169 106
rect -162 103 -160 106
rect 24 92 26 111
rect 34 92 36 111
rect 79 94 81 97
rect 89 94 91 97
rect -195 85 -193 86
rect -189 83 -187 86
rect -112 75 -110 78
rect -106 75 -104 82
rect -90 75 -88 87
rect 24 79 26 82
rect 34 79 36 82
rect -74 75 -72 78
rect -28 71 -26 79
rect 24 71 26 74
rect 34 71 36 74
rect -90 52 -88 55
rect -74 50 -72 55
rect 321 118 323 121
rect 407 115 409 127
rect 447 121 449 133
rect 365 111 367 114
rect 196 107 198 110
rect 325 105 327 108
rect 221 99 223 102
rect 231 99 233 102
rect 162 90 164 93
rect 172 90 174 93
rect 114 74 116 77
rect 138 73 140 77
rect 148 73 150 77
rect -80 39 -78 42
rect -28 44 -26 51
rect -74 39 -72 40
rect -56 39 -54 40
rect -47 39 -45 42
rect -112 23 -110 35
rect -106 32 -104 35
rect -112 10 -110 13
rect -28 37 -26 40
rect 24 31 26 51
rect 34 31 36 51
rect 79 36 81 54
rect 89 36 91 54
rect 114 40 116 54
rect 407 102 409 105
rect 486 112 488 115
rect 492 112 494 119
rect 508 112 510 124
rect 524 112 526 115
rect 447 98 449 101
rect 256 79 258 82
rect 325 73 327 85
rect 365 79 367 91
rect 325 60 327 63
rect 570 108 572 116
rect 508 89 510 92
rect 524 87 526 92
rect 518 76 520 79
rect 570 81 572 88
rect 524 76 526 77
rect 542 76 544 77
rect 551 76 553 79
rect 486 60 488 72
rect 492 69 494 72
rect -28 24 -26 27
rect -56 16 -54 19
rect -47 16 -45 19
rect 138 34 140 53
rect 148 34 150 53
rect 221 41 223 59
rect 231 41 233 59
rect 256 45 258 59
rect 365 56 367 59
rect 486 47 488 50
rect 114 27 116 30
rect 79 23 81 26
rect 89 23 91 26
rect 570 74 572 77
rect 570 61 572 64
rect 542 53 544 56
rect 551 53 553 56
rect 518 35 520 36
rect 256 32 258 35
rect 524 33 526 36
rect 221 28 223 31
rect 231 28 233 31
rect 138 11 140 14
rect 148 11 150 14
rect 24 7 26 11
rect 34 7 36 11
rect -80 -2 -78 -1
rect -74 -4 -72 -1
<< polycontact >>
rect -56 832 -52 836
rect -8 822 -4 826
rect -94 806 -90 810
rect 223 815 227 819
rect 347 819 351 823
rect 395 809 399 813
rect -25 794 -21 798
rect 211 793 215 797
rect 240 796 244 800
rect -60 776 -56 780
rect 309 793 313 797
rect 378 781 382 785
rect 343 763 347 767
rect -56 721 -52 725
rect 61 724 65 728
rect 71 717 75 721
rect 213 725 217 729
rect -8 711 -4 715
rect -94 695 -90 699
rect -169 661 -165 665
rect -25 683 -21 687
rect -60 665 -56 669
rect 326 707 330 711
rect 405 713 409 717
rect 102 692 106 696
rect 314 685 318 689
rect 343 688 347 692
rect 393 691 397 695
rect 422 694 426 698
rect -121 651 -117 655
rect -207 635 -203 639
rect 24 640 28 644
rect 34 647 38 651
rect -138 623 -134 627
rect 505 664 509 668
rect 553 654 557 658
rect -173 605 -169 609
rect -66 582 -62 586
rect 93 604 97 608
rect 103 610 107 614
rect 128 608 132 612
rect 316 617 320 621
rect 395 623 399 627
rect 467 638 471 642
rect 24 585 28 589
rect 34 593 38 597
rect 536 626 540 630
rect 501 608 505 612
rect 159 585 163 589
rect -18 572 -14 576
rect -104 556 -100 560
rect -177 520 -173 524
rect 169 578 173 582
rect -35 544 -31 548
rect -70 526 -66 530
rect -129 510 -125 514
rect -215 494 -211 498
rect -146 482 -142 486
rect 324 535 328 539
rect 415 535 419 539
rect 93 506 97 510
rect 103 512 107 516
rect 312 513 316 517
rect 341 516 345 520
rect 151 500 155 504
rect 161 493 165 497
rect 185 500 189 504
rect -181 464 -177 468
rect 19 466 23 470
rect 29 473 33 477
rect -68 421 -64 425
rect 403 513 407 517
rect 432 516 436 520
rect -20 411 -16 415
rect 19 411 23 415
rect -106 395 -102 399
rect -192 367 -188 371
rect 29 419 33 423
rect 83 416 87 420
rect 93 422 97 426
rect 118 420 122 424
rect 314 445 318 449
rect 517 486 521 490
rect 565 476 569 480
rect 405 445 409 449
rect 479 460 483 464
rect 548 448 552 452
rect 513 430 517 434
rect 206 411 210 415
rect 216 417 220 421
rect 241 415 245 419
rect -37 383 -33 387
rect 156 398 160 402
rect 166 391 170 395
rect -72 365 -68 369
rect -144 357 -140 361
rect -230 341 -226 345
rect -161 329 -157 333
rect -196 311 -192 315
rect 329 369 333 373
rect 416 369 420 373
rect 317 347 321 351
rect 346 350 350 354
rect 74 318 78 322
rect 84 324 88 328
rect 18 293 22 297
rect 28 300 32 304
rect 404 347 408 351
rect 433 350 437 354
rect 195 305 199 309
rect 205 298 209 302
rect 229 305 233 309
rect -75 248 -71 252
rect -27 238 -23 242
rect 18 238 22 242
rect -113 222 -109 226
rect 28 246 32 250
rect 319 279 323 283
rect 517 329 521 333
rect 565 319 569 323
rect 479 303 483 307
rect 406 279 410 283
rect 548 291 552 295
rect 513 273 517 277
rect -44 210 -40 214
rect 81 225 85 229
rect 91 231 95 235
rect 116 229 120 233
rect 156 206 160 210
rect 166 199 170 203
rect -79 192 -75 196
rect -193 137 -189 141
rect -145 127 -141 131
rect -231 111 -227 115
rect 201 194 205 198
rect 211 200 215 204
rect 236 198 240 202
rect 413 206 417 210
rect 517 210 521 214
rect 565 200 569 204
rect 401 184 405 188
rect 430 187 434 191
rect 331 164 335 168
rect 479 184 483 188
rect 548 172 552 176
rect 513 154 517 158
rect 81 127 85 131
rect 91 133 95 137
rect 319 142 323 146
rect 348 145 352 149
rect 158 121 162 125
rect 168 114 172 118
rect 192 121 196 125
rect -162 99 -158 103
rect 20 93 24 97
rect 30 100 34 104
rect -197 81 -193 85
rect -78 50 -74 54
rect 403 116 407 120
rect -30 40 -26 44
rect -116 24 -112 28
rect 20 38 24 42
rect 30 46 34 50
rect 75 37 79 41
rect 85 43 89 47
rect 110 41 114 45
rect 321 74 325 78
rect 520 87 524 91
rect 568 77 572 81
rect 482 61 486 65
rect 134 42 138 46
rect -47 12 -43 16
rect 144 35 148 39
rect 217 42 221 46
rect 227 48 231 52
rect 252 46 256 50
rect 551 49 555 53
rect 516 31 520 35
rect -82 -6 -78 -2
<< polynpluscontact >>
rect 253 731 257 735
rect 356 623 360 627
rect 435 629 439 633
rect 354 451 358 455
rect 445 451 449 455
rect 359 285 363 289
rect 446 285 450 289
rect 443 122 447 126
rect 361 80 365 84
<< metal1 >>
rect -95 872 -8 875
rect -95 857 -91 872
rect -73 857 -69 872
rect -57 857 -53 872
rect -11 853 -8 872
rect 308 859 395 862
rect 201 853 255 856
rect -45 840 -36 841
rect -45 837 -12 840
rect -65 836 -61 837
rect -65 832 -56 836
rect -65 829 -61 832
rect -69 826 -59 829
rect -105 806 -94 810
rect -81 808 -77 817
rect -87 805 -77 808
rect -95 773 -91 795
rect -80 779 -77 805
rect -69 798 -66 826
rect -63 821 -59 826
rect -41 821 -38 837
rect -15 826 -12 837
rect -1 826 3 833
rect -15 823 -8 826
rect -1 822 49 826
rect -1 819 3 822
rect -69 794 -25 798
rect -80 776 -60 779
rect -49 773 -45 781
rect -18 773 -15 801
rect -11 773 -8 809
rect -95 770 -8 773
rect -95 761 -8 764
rect -95 746 -91 761
rect -73 746 -69 761
rect -57 746 -53 761
rect -11 742 -8 761
rect -45 729 -36 730
rect 45 729 49 822
rect 201 777 204 853
rect 222 846 225 853
rect 212 815 223 818
rect 231 818 234 826
rect 231 815 243 818
rect 207 797 210 815
rect 231 814 234 815
rect 222 800 225 804
rect 240 800 243 815
rect 222 797 227 800
rect 207 794 211 797
rect 246 772 249 775
rect 217 769 249 772
rect 60 762 82 765
rect 201 763 217 766
rect 60 755 63 762
rect 79 755 82 762
rect 212 756 215 763
rect -45 726 -12 729
rect -65 725 -61 726
rect -65 721 -56 725
rect -65 718 -61 721
rect -69 715 -59 718
rect -208 701 -121 704
rect -208 686 -204 701
rect -186 686 -182 701
rect -170 686 -166 701
rect -124 682 -121 701
rect -106 695 -94 699
rect -81 697 -77 706
rect -87 694 -77 697
rect -158 669 -149 670
rect -158 666 -125 669
rect -178 665 -174 666
rect -178 661 -169 665
rect -178 658 -174 661
rect -182 655 -172 658
rect -218 635 -207 639
rect -194 637 -190 646
rect -200 634 -190 637
rect -208 602 -204 624
rect -193 608 -190 634
rect -182 627 -179 655
rect -176 650 -172 655
rect -154 650 -151 666
rect -128 655 -125 666
rect -114 655 -110 662
rect -95 662 -91 684
rect -80 668 -77 694
rect -69 687 -66 715
rect -63 710 -59 715
rect -41 710 -38 726
rect -15 715 -12 726
rect 49 724 61 727
rect 70 727 73 735
rect 96 730 106 733
rect 70 724 88 727
rect -1 715 3 722
rect 32 716 42 720
rect 32 715 36 716
rect 47 717 71 720
rect 79 716 82 724
rect -15 712 -8 715
rect -1 711 36 715
rect -1 708 3 711
rect 17 704 46 708
rect 23 698 27 704
rect -69 683 -25 687
rect -80 665 -60 668
rect -49 662 -45 670
rect -18 662 -15 690
rect -11 662 -8 698
rect 60 693 63 696
rect 85 695 88 724
rect 101 723 104 730
rect 206 725 213 728
rect 221 728 224 736
rect 246 734 249 769
rect 252 762 255 853
rect 308 844 312 859
rect 330 844 334 859
rect 346 844 350 859
rect 392 840 395 859
rect 358 827 367 828
rect 358 824 391 827
rect 338 823 342 824
rect 338 819 347 823
rect 338 816 342 819
rect 334 813 344 816
rect 305 796 309 797
rect 289 793 309 796
rect 322 795 326 804
rect 246 731 253 734
rect 261 734 264 742
rect 289 734 292 793
rect 316 792 326 795
rect 308 760 312 782
rect 323 766 326 792
rect 334 785 337 813
rect 340 808 344 813
rect 362 808 365 824
rect 388 813 391 824
rect 402 813 406 820
rect 388 810 395 813
rect 402 809 418 813
rect 402 806 406 809
rect 334 781 378 785
rect 323 763 343 766
rect 354 760 358 768
rect 385 760 388 788
rect 392 760 395 796
rect 308 757 395 760
rect 383 751 437 754
rect 261 731 292 734
rect 304 745 358 748
rect 261 730 264 731
rect 221 725 236 728
rect 221 724 224 725
rect 212 707 215 714
rect 252 707 255 710
rect 212 704 227 707
rect 110 696 113 703
rect 232 704 255 707
rect 59 690 64 693
rect 81 692 102 695
rect 110 693 150 696
rect -95 659 -8 662
rect -128 652 -121 655
rect -114 652 -100 655
rect -114 651 -108 652
rect -114 648 -110 651
rect 8 647 34 651
rect -182 623 -138 627
rect -193 605 -173 608
rect -162 602 -158 610
rect -131 602 -128 630
rect -124 602 -121 638
rect -105 622 -18 625
rect 8 623 11 647
rect 41 644 45 658
rect -105 607 -101 622
rect -83 607 -79 622
rect -67 607 -63 622
rect -21 603 -18 622
rect -208 599 -121 602
rect -55 590 -46 591
rect -55 587 -22 590
rect 8 589 11 618
rect 14 640 24 644
rect 32 640 72 644
rect 32 639 36 640
rect 14 597 17 635
rect 23 625 27 629
rect 41 625 45 629
rect 23 622 45 625
rect 23 618 27 622
rect 68 607 72 640
rect 85 614 88 692
rect 110 691 113 693
rect 101 677 104 681
rect 101 674 111 677
rect 92 668 125 671
rect 304 669 307 745
rect 325 738 328 745
rect 315 707 326 710
rect 334 710 337 718
rect 334 707 346 710
rect 310 689 313 707
rect 334 706 337 707
rect 325 692 328 696
rect 343 692 346 707
rect 325 689 330 692
rect 310 686 314 689
rect 92 661 95 668
rect 122 651 125 668
rect 349 664 352 667
rect 320 661 352 664
rect 304 655 320 658
rect 122 648 130 651
rect 127 641 130 648
rect 315 648 318 655
rect 85 611 103 614
rect 111 612 114 621
rect 136 612 139 621
rect 158 623 180 626
rect 158 616 161 623
rect 177 616 180 623
rect 309 617 316 620
rect 324 620 327 628
rect 349 626 352 661
rect 355 654 358 745
rect 383 675 386 751
rect 404 744 407 751
rect 389 713 405 716
rect 413 716 416 724
rect 413 713 425 716
rect 389 704 392 713
rect 413 712 416 713
rect 389 695 392 699
rect 404 698 407 702
rect 422 698 425 713
rect 404 695 409 698
rect 389 692 393 695
rect 428 670 431 673
rect 399 667 431 670
rect 383 661 399 664
rect 394 654 397 661
rect 349 623 356 626
rect 364 626 367 634
rect 364 623 383 626
rect 364 622 367 623
rect 324 617 339 620
rect 388 623 395 626
rect 403 626 406 634
rect 428 632 431 667
rect 434 660 437 751
rect 466 704 553 707
rect 466 689 470 704
rect 488 689 492 704
rect 504 689 508 704
rect 550 685 553 704
rect 516 672 525 673
rect 516 669 549 672
rect 496 668 500 669
rect 496 664 505 668
rect 496 661 500 664
rect 492 658 502 661
rect 428 629 435 632
rect 443 632 446 640
rect 459 638 467 642
rect 480 640 484 649
rect 459 632 462 638
rect 474 637 484 640
rect 443 629 462 632
rect 443 628 446 629
rect 403 623 418 626
rect 403 622 406 623
rect 324 616 327 617
rect 111 609 128 612
rect 68 604 78 607
rect 83 604 93 607
rect 111 607 114 609
rect 136 609 145 612
rect 136 607 139 609
rect 102 604 114 607
rect 102 603 105 604
rect 14 593 34 597
rect 41 589 45 598
rect -75 586 -71 587
rect -75 582 -66 586
rect -75 579 -71 582
rect -79 576 -69 579
rect -216 560 -129 563
rect -216 545 -212 560
rect -194 545 -190 560
rect -178 545 -174 560
rect -132 541 -129 560
rect -118 556 -104 560
rect -91 558 -87 567
rect -97 555 -87 558
rect -166 528 -157 529
rect -166 525 -133 528
rect -186 524 -182 525
rect -186 520 -177 524
rect -186 517 -182 520
rect -190 514 -180 517
rect -219 497 -215 498
rect -226 494 -215 497
rect -202 496 -198 505
rect -208 493 -198 496
rect -216 461 -212 483
rect -201 467 -198 493
rect -190 486 -187 514
rect -184 509 -180 514
rect -162 509 -159 525
rect -136 514 -133 525
rect -122 514 -118 521
rect -105 523 -101 545
rect -90 529 -87 555
rect -79 548 -76 576
rect -73 571 -69 576
rect -51 571 -48 587
rect -25 576 -22 587
rect -11 576 -7 583
rect 8 585 24 589
rect 32 585 67 589
rect 8 576 11 585
rect -25 573 -18 576
rect -11 572 11 576
rect 32 578 36 585
rect 63 581 67 585
rect 92 587 95 593
rect 111 587 114 593
rect 127 587 130 597
rect 92 584 130 587
rect 142 588 145 609
rect 315 599 318 606
rect 394 605 397 612
rect 434 605 437 608
rect 394 602 409 605
rect 355 599 358 602
rect 414 602 437 605
rect 466 605 470 627
rect 481 611 484 637
rect 492 630 495 658
rect 498 653 502 658
rect 520 653 523 669
rect 546 658 549 669
rect 560 658 564 665
rect 546 655 553 658
rect 560 654 574 658
rect 560 651 564 654
rect 492 626 536 630
rect 481 608 501 611
rect 512 605 516 613
rect 543 605 546 633
rect 550 605 553 641
rect 466 602 553 605
rect 315 596 330 599
rect 142 585 159 588
rect 168 588 171 596
rect 335 596 358 599
rect 168 585 189 588
rect 60 578 169 581
rect 177 577 180 585
rect 90 572 96 575
rect 302 573 356 576
rect -11 569 -7 572
rect 92 563 95 572
rect -79 544 -35 548
rect -90 526 -70 529
rect -59 523 -55 531
rect -28 523 -25 551
rect -21 523 -18 559
rect 23 550 27 558
rect 41 552 45 558
rect 158 554 161 557
rect 41 550 46 552
rect 23 547 46 550
rect 157 551 162 554
rect 150 538 187 541
rect 12 530 41 534
rect 150 531 153 538
rect 169 531 172 538
rect -105 520 -18 523
rect 18 524 22 530
rect 184 531 187 538
rect -136 511 -129 514
rect -122 513 -116 514
rect 84 513 103 516
rect -122 510 -103 513
rect -122 507 -118 510
rect 111 514 114 523
rect 111 511 122 514
rect 48 506 64 509
rect 69 506 93 509
rect 111 509 114 511
rect 102 506 114 509
rect -190 482 -146 486
rect -201 464 -181 467
rect -170 461 -166 469
rect -139 461 -136 489
rect -132 461 -129 497
rect 3 473 29 477
rect -216 458 -129 461
rect -107 461 -20 464
rect -107 446 -103 461
rect -85 446 -81 461
rect -69 446 -65 461
rect -23 442 -20 461
rect 3 450 6 473
rect 36 470 40 484
rect 48 470 51 506
rect -57 429 -48 430
rect -57 426 -24 429
rect -77 425 -73 426
rect -77 421 -68 425
rect -77 418 -73 421
rect -81 415 -71 418
rect -231 407 -144 410
rect -231 392 -227 407
rect -209 392 -205 407
rect -193 392 -189 407
rect -147 388 -144 407
rect -122 395 -106 399
rect -93 397 -89 406
rect -99 394 -89 397
rect -181 375 -172 376
rect -181 372 -148 375
rect -201 371 -197 372
rect -201 367 -192 371
rect -201 364 -197 367
rect -205 361 -195 364
rect -242 341 -230 345
rect -217 343 -213 352
rect -223 340 -213 343
rect -231 308 -227 330
rect -216 314 -213 340
rect -205 333 -202 361
rect -199 356 -195 361
rect -177 356 -174 372
rect -151 361 -148 372
rect -137 361 -133 368
rect -107 362 -103 384
rect -92 368 -89 394
rect -81 387 -78 415
rect -75 410 -71 415
rect -53 410 -50 426
rect -27 415 -24 426
rect -13 415 -9 422
rect 3 415 6 445
rect 14 466 19 470
rect 27 466 51 470
rect 27 465 31 466
rect 9 423 12 465
rect 18 451 22 455
rect 36 451 40 455
rect 18 448 40 451
rect 18 444 22 448
rect 9 419 29 423
rect 36 415 40 424
rect 75 426 78 506
rect 102 505 105 506
rect 92 489 95 495
rect 111 489 114 495
rect 119 496 122 511
rect 140 500 151 503
rect 160 503 163 511
rect 193 504 196 511
rect 160 500 185 503
rect 193 501 202 504
rect 119 493 161 496
rect 169 492 172 500
rect 193 499 196 501
rect 92 486 114 489
rect 82 480 115 483
rect 82 473 85 480
rect 112 463 115 480
rect 150 469 153 472
rect 184 469 187 489
rect 149 466 187 469
rect 112 460 120 463
rect 117 453 120 460
rect 75 423 93 426
rect 101 424 104 433
rect 126 424 129 433
rect 155 436 177 439
rect 155 429 158 436
rect 174 429 177 436
rect 101 421 118 424
rect 62 416 83 419
rect 101 419 104 421
rect 126 421 135 424
rect 199 421 202 501
rect 302 497 305 573
rect 323 566 326 573
rect 313 535 324 538
rect 332 538 335 546
rect 332 535 344 538
rect 308 517 311 535
rect 332 534 335 535
rect 323 520 326 524
rect 341 520 344 535
rect 323 517 328 520
rect 308 514 312 517
rect 347 492 350 495
rect 318 489 350 492
rect 302 483 318 486
rect 205 475 238 478
rect 205 468 208 475
rect 235 458 238 475
rect 313 476 316 483
rect 235 455 243 458
rect 240 448 243 455
rect 307 445 314 448
rect 322 448 325 456
rect 347 454 350 489
rect 353 482 356 573
rect 393 573 447 576
rect 393 497 396 573
rect 414 566 417 573
rect 404 535 415 538
rect 423 538 426 546
rect 423 535 435 538
rect 399 517 402 535
rect 423 534 426 535
rect 414 520 417 524
rect 432 520 435 535
rect 414 517 419 520
rect 399 514 403 517
rect 438 492 441 495
rect 409 489 441 492
rect 393 483 409 486
rect 404 476 407 483
rect 347 451 354 454
rect 362 454 365 462
rect 362 451 371 454
rect 362 450 365 451
rect 322 445 337 448
rect 368 448 371 451
rect 368 445 393 448
rect 322 444 325 445
rect 398 445 405 448
rect 413 448 416 456
rect 438 454 441 489
rect 444 482 447 573
rect 478 526 565 529
rect 478 511 482 526
rect 500 511 504 526
rect 516 511 520 526
rect 562 507 565 526
rect 528 494 537 495
rect 528 491 561 494
rect 508 490 512 491
rect 508 486 517 490
rect 508 483 512 486
rect 504 480 514 483
rect 438 451 445 454
rect 453 454 456 462
rect 469 460 479 464
rect 492 462 496 471
rect 469 454 472 460
rect 486 459 496 462
rect 453 451 472 454
rect 453 450 456 451
rect 413 445 428 448
rect 413 444 416 445
rect 126 419 129 421
rect 92 416 104 419
rect 92 415 95 416
rect -27 412 -20 415
rect -13 411 19 415
rect 27 411 52 415
rect -13 408 -9 411
rect 27 404 31 411
rect -81 383 -37 387
rect -92 365 -72 368
rect -61 362 -57 370
rect -30 362 -27 390
rect -23 362 -20 398
rect 49 393 52 411
rect 82 399 85 405
rect 101 399 104 405
rect 117 399 120 409
rect 82 396 120 399
rect 132 401 135 421
rect 198 418 216 421
rect 224 419 227 428
rect 249 419 252 428
rect 313 427 316 434
rect 353 427 356 430
rect 313 424 328 427
rect 333 424 356 427
rect 404 427 407 434
rect 444 427 447 430
rect 404 424 419 427
rect 424 424 447 427
rect 478 427 482 449
rect 493 433 496 459
rect 504 452 507 480
rect 510 475 514 480
rect 532 475 535 491
rect 558 480 561 491
rect 572 480 576 487
rect 558 477 565 480
rect 572 476 585 480
rect 572 473 576 476
rect 504 448 548 452
rect 493 430 513 433
rect 524 427 528 435
rect 555 427 558 455
rect 562 427 565 463
rect 478 424 565 427
rect 224 416 241 419
rect 132 398 156 401
rect 165 401 168 409
rect 194 411 206 414
rect 224 414 227 416
rect 249 416 258 419
rect 249 414 252 416
rect 215 411 227 414
rect 194 401 197 411
rect 215 410 218 411
rect 307 407 361 410
rect 165 398 197 401
rect 49 390 73 393
rect 148 393 166 394
rect 78 391 166 393
rect 78 390 151 391
rect 174 390 177 398
rect 205 394 208 400
rect 224 394 227 400
rect 240 394 243 404
rect 205 391 243 394
rect 18 376 22 384
rect 71 384 77 387
rect 36 378 40 384
rect 36 376 41 378
rect 18 373 41 376
rect 73 375 76 384
rect 155 367 158 370
rect 154 364 159 367
rect -151 358 -144 361
rect -137 360 -131 361
rect -137 357 -119 360
rect -107 359 -20 362
rect 11 357 40 361
rect -137 354 -133 357
rect 17 351 21 357
rect -205 329 -161 333
rect -216 311 -196 314
rect -185 308 -181 316
rect -154 308 -151 336
rect -147 308 -144 344
rect 194 343 231 346
rect 65 325 84 328
rect 92 326 95 335
rect 194 336 197 343
rect 213 336 216 343
rect 228 336 231 343
rect 307 331 310 407
rect 328 400 331 407
rect 318 369 329 372
rect 337 372 340 380
rect 337 369 349 372
rect 313 351 316 369
rect 337 368 340 369
rect 328 354 331 358
rect 346 354 349 369
rect 328 351 333 354
rect 313 348 317 351
rect 352 326 355 329
rect 92 323 145 326
rect 323 323 355 326
rect 48 318 74 321
rect 92 321 95 323
rect 83 318 95 321
rect -231 305 -144 308
rect 2 300 28 304
rect -114 288 -27 291
rect -114 273 -110 288
rect -92 273 -88 288
rect -76 273 -72 288
rect -30 269 -27 288
rect 2 284 5 300
rect 35 297 39 311
rect 48 297 52 318
rect -64 256 -55 257
rect -64 253 -31 256
rect -84 252 -80 253
rect -84 248 -75 252
rect -84 245 -80 248
rect -88 242 -78 245
rect -130 222 -113 226
rect -100 224 -96 233
rect -106 221 -96 224
rect -114 189 -110 211
rect -99 195 -96 221
rect -88 214 -85 242
rect -82 237 -78 242
rect -60 237 -57 253
rect -34 242 -31 253
rect -20 242 -16 249
rect 2 242 5 279
rect 13 293 18 297
rect 26 293 52 297
rect 26 292 30 293
rect 8 250 11 292
rect 17 278 21 282
rect 35 278 39 282
rect 17 275 39 278
rect 17 271 21 275
rect 8 246 28 250
rect 35 242 39 251
rect -34 239 -27 242
rect -20 238 18 242
rect 26 238 49 242
rect -20 235 -16 238
rect 26 231 30 238
rect 61 228 64 318
rect 83 317 86 318
rect 73 301 76 307
rect 92 301 95 307
rect 73 298 95 301
rect 142 301 145 323
rect 307 317 323 320
rect 186 305 195 308
rect 204 308 207 316
rect 237 309 240 316
rect 318 310 321 317
rect 204 305 229 308
rect 237 306 246 309
rect 142 298 205 301
rect 213 297 216 305
rect 237 304 240 306
rect 80 289 113 292
rect 80 282 83 289
rect 110 272 113 289
rect 194 274 197 277
rect 228 274 231 294
rect 110 269 118 272
rect 193 271 231 274
rect 115 262 118 269
rect 243 268 246 306
rect 312 279 319 282
rect 327 282 330 290
rect 352 288 355 323
rect 358 316 361 407
rect 394 407 448 410
rect 394 331 397 407
rect 415 400 418 407
rect 405 369 416 372
rect 424 372 427 380
rect 424 369 436 372
rect 400 351 403 369
rect 424 368 427 369
rect 415 354 418 358
rect 433 354 436 369
rect 415 351 420 354
rect 400 348 404 351
rect 439 326 442 329
rect 410 323 442 326
rect 394 317 410 320
rect 405 310 408 317
rect 352 285 359 288
rect 367 288 370 296
rect 367 285 389 288
rect 367 284 370 285
rect 327 279 342 282
rect 386 282 389 285
rect 386 279 394 282
rect 327 278 330 279
rect 399 279 406 282
rect 414 282 417 290
rect 439 288 442 323
rect 445 316 448 407
rect 478 369 565 372
rect 478 354 482 369
rect 500 354 504 369
rect 516 354 520 369
rect 562 350 565 369
rect 528 337 537 338
rect 528 334 561 337
rect 508 333 512 334
rect 508 329 517 333
rect 508 326 512 329
rect 504 323 514 326
rect 471 303 479 307
rect 492 305 496 314
rect 439 285 446 288
rect 454 288 457 296
rect 471 288 474 303
rect 486 302 496 305
rect 454 285 474 288
rect 454 284 457 285
rect 414 279 429 282
rect 414 278 417 279
rect 194 265 246 268
rect 478 270 482 292
rect 493 276 496 302
rect 504 295 507 323
rect 510 318 514 323
rect 532 318 535 334
rect 558 323 561 334
rect 572 323 576 330
rect 558 320 565 323
rect 572 319 587 323
rect 572 316 576 319
rect 504 291 548 295
rect 493 273 513 276
rect 524 270 528 278
rect 555 270 558 298
rect 562 270 565 306
rect 72 232 91 235
rect 99 233 102 242
rect 124 233 127 242
rect 155 244 177 247
rect 155 237 158 244
rect 174 237 177 244
rect 99 230 116 233
rect 61 225 81 228
rect 99 228 102 230
rect 124 230 133 233
rect 124 228 127 230
rect 90 225 102 228
rect -88 210 -44 214
rect -99 192 -79 195
rect -68 189 -64 197
rect -37 189 -34 217
rect -30 189 -27 225
rect 17 203 21 211
rect 35 205 39 211
rect 35 203 40 205
rect 17 200 40 203
rect -114 186 -27 189
rect -232 177 -145 180
rect -232 162 -228 177
rect -210 162 -206 177
rect -194 162 -190 177
rect -148 158 -145 177
rect 13 157 42 161
rect 19 151 23 157
rect -182 145 -173 146
rect -182 142 -149 145
rect -202 141 -198 142
rect -202 137 -193 141
rect -202 134 -198 137
rect -206 131 -196 134
rect -248 111 -231 115
rect -218 113 -214 122
rect -224 110 -214 113
rect -232 78 -228 100
rect -217 84 -214 110
rect -206 103 -203 131
rect -200 126 -196 131
rect -178 126 -175 142
rect -152 131 -149 142
rect -138 131 -134 138
rect 61 137 64 225
rect 90 224 93 225
rect 80 208 83 214
rect 99 208 102 214
rect 115 208 118 218
rect 80 205 118 208
rect 130 209 133 230
rect 130 206 156 209
rect 165 209 168 217
rect 165 206 183 209
rect 73 199 166 202
rect 174 198 177 206
rect 78 193 84 196
rect 180 197 183 206
rect 194 204 197 265
rect 318 261 321 268
rect 358 261 361 264
rect 200 258 233 261
rect 318 258 333 261
rect 200 251 203 258
rect 230 241 233 258
rect 338 258 361 261
rect 405 261 408 268
rect 478 267 565 270
rect 445 261 448 264
rect 405 258 420 261
rect 425 258 448 261
rect 478 250 565 253
rect 391 244 445 247
rect 230 238 238 241
rect 235 231 238 238
rect 194 201 211 204
rect 219 202 222 211
rect 244 202 247 211
rect 219 199 236 202
rect 180 194 201 197
rect 219 197 222 199
rect 244 199 251 202
rect 309 202 363 205
rect 244 197 247 199
rect 210 194 222 197
rect 210 193 213 194
rect 80 184 83 193
rect 155 175 158 178
rect 200 177 203 183
rect 219 177 222 183
rect 235 177 238 187
rect 154 172 159 175
rect 200 174 238 177
rect 157 159 194 162
rect 157 152 160 159
rect 176 152 179 159
rect 191 152 194 159
rect 61 134 91 137
rect 99 135 102 144
rect 99 132 134 135
rect -152 128 -145 131
rect -138 127 -123 131
rect 61 127 81 130
rect 99 130 102 132
rect 90 127 102 130
rect -138 124 -134 127
rect -206 99 -162 103
rect -217 81 -197 84
rect -186 78 -182 86
rect -155 78 -152 106
rect -148 78 -145 114
rect 4 100 30 104
rect -232 75 -145 78
rect -117 90 -30 93
rect -117 75 -113 90
rect -95 75 -91 90
rect -79 75 -75 90
rect -33 71 -30 90
rect 4 79 7 100
rect 37 97 41 111
rect 61 97 64 127
rect 90 126 93 127
rect 80 110 83 116
rect 99 110 102 116
rect 131 117 134 132
rect 150 121 158 124
rect 167 124 170 132
rect 200 125 203 132
rect 309 126 312 202
rect 330 195 333 202
rect 320 164 331 167
rect 339 167 342 175
rect 339 164 351 167
rect 339 163 342 164
rect 315 146 318 162
rect 330 149 333 153
rect 348 149 351 164
rect 330 146 335 149
rect 315 143 319 146
rect 167 121 192 124
rect 200 122 209 125
rect 131 114 168 117
rect 176 113 179 121
rect 200 120 203 122
rect 80 107 102 110
rect -67 58 -58 59
rect -67 55 -34 58
rect -87 54 -83 55
rect -87 50 -78 54
rect -87 47 -83 50
rect -91 44 -81 47
rect -136 24 -116 28
rect -103 26 -99 35
rect -109 23 -99 26
rect -117 -9 -113 13
rect -102 -3 -99 23
rect -91 16 -88 44
rect -85 39 -81 44
rect -63 39 -60 55
rect -37 44 -34 55
rect -23 44 -19 51
rect 4 44 7 74
rect 15 93 20 97
rect 28 93 64 97
rect 28 92 32 93
rect 10 50 13 92
rect 19 78 23 82
rect 37 78 41 82
rect 19 75 41 78
rect 19 71 23 75
rect 61 63 64 93
rect 74 101 107 104
rect 74 94 77 101
rect 104 84 107 101
rect 157 90 160 93
rect 191 90 194 110
rect 156 87 194 90
rect 104 81 112 84
rect 109 74 112 81
rect 133 80 155 83
rect 133 73 136 80
rect 152 73 155 80
rect 53 60 64 63
rect 10 46 30 50
rect -37 41 -30 44
rect -23 42 7 44
rect 37 42 41 51
rect -23 40 20 42
rect -23 37 -19 40
rect 4 38 20 40
rect 28 38 47 42
rect 28 31 32 38
rect -91 12 -47 16
rect -102 -6 -82 -3
rect -71 -9 -67 -1
rect -40 -9 -37 19
rect -33 -9 -30 27
rect 19 3 23 11
rect 37 5 41 11
rect 44 11 47 38
rect 53 40 56 60
rect 65 44 85 47
rect 93 45 96 54
rect 118 45 121 54
rect 93 42 110 45
rect 53 37 75 40
rect 93 40 96 42
rect 118 42 134 45
rect 143 45 146 53
rect 206 52 209 122
rect 354 121 357 124
rect 325 118 357 121
rect 309 112 325 115
rect 216 106 249 109
rect 216 99 219 106
rect 246 89 249 106
rect 320 105 323 112
rect 246 86 254 89
rect 251 79 254 86
rect 314 74 321 77
rect 329 77 332 85
rect 354 83 357 118
rect 360 111 363 202
rect 391 168 394 244
rect 412 237 415 244
rect 397 206 413 209
rect 421 209 424 217
rect 421 206 433 209
rect 397 203 400 206
rect 421 205 424 206
rect 397 188 400 198
rect 412 191 415 195
rect 430 191 433 206
rect 412 188 417 191
rect 397 185 401 188
rect 436 163 439 166
rect 407 160 439 163
rect 391 154 407 157
rect 402 147 405 154
rect 396 116 403 119
rect 411 119 414 127
rect 436 125 439 160
rect 442 153 445 244
rect 478 235 482 250
rect 500 235 504 250
rect 516 235 520 250
rect 562 231 565 250
rect 528 218 537 219
rect 528 215 561 218
rect 508 214 512 215
rect 508 210 517 214
rect 508 207 512 210
rect 504 204 514 207
rect 469 185 479 188
rect 436 122 443 125
rect 451 125 454 133
rect 469 125 472 185
rect 475 184 479 185
rect 492 186 496 195
rect 486 183 496 186
rect 478 151 482 173
rect 493 157 496 183
rect 504 176 507 204
rect 510 199 514 204
rect 532 199 535 215
rect 558 204 561 215
rect 572 204 576 211
rect 558 201 565 204
rect 572 200 589 204
rect 572 197 576 200
rect 504 172 548 176
rect 493 154 513 157
rect 524 151 528 159
rect 555 151 558 179
rect 562 151 565 187
rect 478 148 565 151
rect 451 122 472 125
rect 481 127 568 130
rect 451 121 454 122
rect 411 116 426 119
rect 411 115 414 116
rect 354 80 361 83
rect 369 83 372 91
rect 391 83 394 114
rect 481 112 485 127
rect 503 112 507 127
rect 519 112 523 127
rect 565 108 568 127
rect 402 98 405 105
rect 442 98 445 101
rect 402 95 417 98
rect 422 95 445 98
rect 531 95 540 96
rect 531 92 564 95
rect 511 91 515 92
rect 511 87 520 91
rect 511 84 515 87
rect 369 80 394 83
rect 507 81 517 84
rect 369 79 372 80
rect 329 74 344 77
rect 329 73 332 74
rect 206 49 227 52
rect 235 50 238 59
rect 260 50 263 59
rect 320 56 323 63
rect 473 61 482 65
rect 495 63 499 72
rect 360 56 363 59
rect 320 53 335 56
rect 340 53 363 56
rect 235 47 252 50
rect 143 42 217 45
rect 235 45 238 47
rect 260 47 271 50
rect 260 45 263 47
rect 226 42 238 45
rect 118 40 121 42
rect 84 37 96 40
rect 84 36 87 37
rect 124 35 144 38
rect 74 20 77 26
rect 93 20 96 26
rect 109 20 112 30
rect 74 17 112 20
rect 124 11 127 35
rect 152 34 155 42
rect 226 41 229 42
rect 268 43 271 47
rect 473 43 476 61
rect 489 60 499 63
rect 268 40 476 43
rect 216 25 219 31
rect 235 25 238 31
rect 251 25 254 35
rect 481 28 485 50
rect 496 34 499 60
rect 507 53 510 81
rect 513 76 517 81
rect 535 76 538 92
rect 561 81 564 92
rect 575 81 579 88
rect 561 78 568 81
rect 575 77 594 81
rect 575 74 579 77
rect 507 49 551 53
rect 496 31 516 34
rect 527 28 531 36
rect 558 28 561 56
rect 565 28 568 64
rect 481 25 568 28
rect 216 22 254 25
rect 133 11 136 14
rect 44 8 127 11
rect 132 8 137 11
rect 37 3 42 5
rect 19 0 42 3
rect -117 -12 -30 -9
<< m2contact >>
rect 227 795 232 800
rect 46 704 51 709
rect 236 725 241 730
rect 227 702 232 707
rect 150 693 155 698
rect -100 650 -95 655
rect 330 687 335 692
rect 389 699 394 704
rect 409 693 414 698
rect 339 617 344 622
rect 383 621 388 626
rect 418 623 423 628
rect 78 602 83 607
rect 409 600 414 605
rect 330 594 335 599
rect 189 585 194 590
rect 55 576 60 581
rect 46 547 51 552
rect 41 530 46 535
rect 79 513 84 518
rect -103 508 -98 513
rect 64 506 69 511
rect 57 416 62 421
rect 328 515 333 520
rect 399 535 404 540
rect 419 515 424 520
rect 337 445 342 450
rect 393 443 398 448
rect 428 445 433 450
rect 328 422 333 427
rect 419 422 424 427
rect 258 416 263 421
rect 73 390 78 395
rect 41 373 46 378
rect 40 357 45 362
rect -122 352 -117 357
rect 60 325 65 330
rect 333 349 338 354
rect 49 238 54 243
rect 181 305 186 310
rect 400 369 405 374
rect 420 349 425 354
rect 342 279 347 284
rect 394 277 399 282
rect 429 279 434 284
rect 67 232 72 237
rect 40 200 45 205
rect 42 157 47 162
rect 67 199 73 205
rect 333 256 338 261
rect 420 256 425 261
rect -123 127 -118 132
rect 145 121 150 126
rect 335 144 340 149
rect 60 44 65 49
rect 417 186 422 191
rect 391 114 396 119
rect 426 116 431 121
rect 417 93 422 98
rect 344 74 349 79
rect 335 51 340 56
rect 42 0 47 5
<< pm12contact >>
rect -84 864 -79 869
rect -66 864 -61 869
rect -52 822 -47 827
rect -34 822 -29 827
rect -84 753 -79 758
rect -66 753 -61 758
rect -197 693 -192 698
rect -179 693 -174 698
rect -165 651 -160 656
rect -147 651 -142 656
rect -52 711 -47 716
rect -34 711 -29 716
rect 319 851 324 856
rect 337 851 342 856
rect 351 809 356 814
rect 369 809 374 814
rect -94 614 -89 619
rect -76 614 -71 619
rect 477 696 482 701
rect 495 696 500 701
rect -205 552 -200 557
rect -187 552 -182 557
rect -173 510 -168 515
rect -155 510 -150 515
rect -62 572 -57 577
rect -44 572 -39 577
rect 509 654 514 659
rect 527 654 532 659
rect -96 453 -91 458
rect -78 453 -73 458
rect -220 399 -215 404
rect -202 399 -197 404
rect -188 357 -183 362
rect -170 357 -165 362
rect -64 411 -59 416
rect -46 411 -41 416
rect 489 518 494 523
rect 507 518 512 523
rect 521 476 526 481
rect 539 476 544 481
rect -103 280 -98 285
rect -85 280 -80 285
rect -71 238 -66 243
rect -53 238 -48 243
rect 489 361 494 366
rect 507 361 512 366
rect 521 319 526 324
rect 539 319 544 324
rect -221 169 -216 174
rect -203 169 -198 174
rect -189 127 -184 132
rect -171 127 -166 132
rect -106 82 -101 87
rect -88 82 -83 87
rect -74 40 -69 45
rect -56 40 -51 45
rect 489 242 494 247
rect 507 242 512 247
rect 521 200 526 205
rect 539 200 544 205
rect 492 119 497 124
rect 510 119 515 124
rect 524 77 529 82
rect 542 77 547 82
<< psm12contact >>
rect 135 500 140 505
<< ndm12contact >>
rect 207 772 212 777
rect 236 775 241 780
rect 310 664 315 669
rect 339 667 344 672
rect 389 670 394 675
rect 418 673 423 678
rect 308 492 313 497
rect 337 495 342 500
rect 399 492 404 497
rect 428 495 433 500
rect 313 326 318 331
rect 342 329 347 334
rect 400 326 405 331
rect 429 329 434 334
rect 315 121 320 126
rect 344 124 349 129
rect 397 163 402 168
rect 426 166 431 171
<< metal2 >>
rect -79 864 -66 867
rect -76 825 -73 864
rect 324 851 337 854
rect -76 822 -52 825
rect -47 822 -34 825
rect 327 812 330 851
rect 327 809 351 812
rect 356 809 369 812
rect 201 772 207 777
rect -79 753 -66 756
rect -76 714 -73 753
rect 201 728 204 772
rect -76 711 -52 714
rect -47 711 -34 714
rect 229 707 232 795
rect 236 730 239 775
rect -192 693 -179 696
rect -189 654 -186 693
rect -189 651 -165 654
rect -160 651 -147 654
rect -98 640 -95 650
rect -98 637 14 640
rect -89 614 -76 617
rect -86 575 -83 614
rect -86 572 -62 575
rect -57 572 -44 575
rect -200 552 -187 555
rect 48 552 51 704
rect 280 699 389 702
rect 280 696 283 699
rect 155 693 283 696
rect 482 696 495 699
rect -197 513 -194 552
rect -197 510 -173 513
rect -168 510 -155 513
rect -101 469 -98 508
rect -101 466 9 469
rect -91 453 -78 456
rect -88 414 -85 453
rect -88 411 -64 414
rect -59 411 -46 414
rect -215 399 -202 402
rect -212 360 -209 399
rect 43 378 46 530
rect 57 421 60 576
rect 80 518 83 602
rect 150 515 153 693
rect 304 664 310 669
rect 304 620 307 664
rect 332 599 335 687
rect 383 670 389 675
rect 339 622 342 667
rect 383 626 386 670
rect 411 605 414 693
rect 418 628 421 673
rect 485 657 488 696
rect 485 654 509 657
rect 514 654 527 657
rect 135 512 153 515
rect 191 563 194 585
rect 191 560 402 563
rect -212 357 -188 360
rect -183 357 -170 360
rect -122 296 -119 352
rect -122 293 8 296
rect -98 280 -85 283
rect -95 241 -92 280
rect -95 238 -71 241
rect -66 238 -53 241
rect 42 205 45 357
rect 66 335 69 506
rect 135 505 138 512
rect 60 332 69 335
rect 60 330 66 332
rect 75 240 78 390
rect 191 317 194 560
rect 399 540 402 560
rect 494 518 507 521
rect 302 492 308 497
rect 302 448 305 492
rect 330 427 333 515
rect 337 450 340 495
rect 393 492 399 497
rect 393 448 396 492
rect 421 427 424 515
rect 428 450 431 495
rect 497 479 500 518
rect 497 476 521 479
rect 526 476 539 479
rect 183 314 194 317
rect 260 387 263 416
rect 260 384 403 387
rect 183 310 186 314
rect 51 202 54 238
rect 67 237 78 240
rect 51 199 67 202
rect -216 169 -203 172
rect -213 130 -210 169
rect -213 127 -189 130
rect -184 127 -171 130
rect -121 97 -118 127
rect -121 94 10 97
rect -101 82 -88 85
rect -98 43 -95 82
rect -98 40 -74 43
rect -69 40 -56 43
rect 44 5 47 157
rect 67 59 70 199
rect 260 168 263 384
rect 400 374 403 384
rect 494 361 507 364
rect 307 326 313 331
rect 307 282 310 326
rect 335 261 338 349
rect 342 284 345 329
rect 394 326 400 331
rect 394 282 397 326
rect 422 261 425 349
rect 429 284 432 329
rect 497 322 500 361
rect 497 319 521 322
rect 526 319 539 322
rect 494 242 507 245
rect 497 203 500 242
rect 497 200 521 203
rect 526 200 539 203
rect 145 165 263 168
rect 145 126 148 165
rect 391 163 397 168
rect 309 121 315 126
rect 309 77 312 121
rect 62 56 70 59
rect 337 56 340 144
rect 344 79 347 124
rect 391 119 394 163
rect 419 98 422 186
rect 426 121 429 166
rect 497 119 510 122
rect 500 80 503 119
rect 500 77 524 80
rect 529 77 542 80
rect 62 49 65 56
<< m123contact >>
rect 207 815 212 820
rect 44 724 49 729
rect 201 723 206 728
rect 42 715 47 720
rect 310 707 315 712
rect 14 635 19 640
rect 6 618 11 623
rect 9 465 14 470
rect 1 445 6 450
rect 304 615 309 620
rect 8 292 13 297
rect 0 279 5 284
rect 308 535 313 540
rect 302 443 307 448
rect 251 199 256 204
rect 10 92 15 97
rect 2 74 7 79
rect 313 369 318 374
rect 307 277 312 282
rect 397 198 402 203
rect 315 162 320 167
rect 309 72 314 77
<< metal3 >>
rect 193 815 207 820
rect 193 729 197 815
rect 49 724 197 729
rect 201 720 206 723
rect 47 715 206 720
rect 296 707 310 711
rect 296 640 300 707
rect 19 636 300 640
rect 11 619 300 622
rect 11 618 304 619
rect 296 615 304 618
rect 288 535 308 538
rect 288 470 291 535
rect 14 467 291 470
rect 6 445 302 448
rect 292 370 313 373
rect 292 297 295 370
rect 13 294 295 297
rect 5 279 307 282
rect 256 199 397 202
rect 299 162 315 165
rect 299 97 302 162
rect 15 94 302 97
rect 7 74 309 77
<< labels >>
rlabel metal1 100 732 100 732 4 vdd
rlabel metal1 107 675 107 675 1 gnd
rlabel metal1 116 694 116 694 7 c1
rlabel metal1 102 585 102 585 1 gnd
rlabel metal1 107 669 107 669 5 vdd
rlabel metal1 82 693 82 693 3 g0_bar
rlabel metal1 69 605 69 605 3 p1_bar
rlabel metal1 169 624 169 624 5 vdd
rlabel metal1 160 552 160 552 1 gnd
rlabel metal1 69 579 69 579 3 g1_bar
rlabel metal1 183 587 183 587 7 c2
rlabel metal1 93 574 93 574 5 vdd
rlabel metal1 102 487 102 487 1 gnd
rlabel metal1 56 507 56 507 3 p2_bar
rlabel metal1 92 397 92 397 1 gnd
rlabel metal1 97 481 97 481 5 vdd
rlabel metal1 165 540 165 540 1 vdd
rlabel metal1 170 467 170 467 1 gnd
rlabel metal1 157 365 157 365 1 gnd
rlabel metal1 166 437 166 437 5 vdd
rlabel metal1 220 477 220 477 1 vdd
rlabel metal1 221 392 221 392 1 gnd
rlabel metal1 73 385 73 385 1 vdd
rlabel metal1 82 299 82 299 1 gnd
rlabel metal1 93 290 93 290 1 vdd
rlabel metal1 98 206 98 206 1 gnd
rlabel metal1 165 245 165 245 1 vdd
rlabel metal1 157 173 157 173 1 gnd
rlabel metal1 255 417 255 417 7 c3
rlabel metal1 209 345 209 345 1 vdd
rlabel metal1 214 273 214 273 1 gnd
rlabel metal1 219 175 219 175 1 gnd
rlabel metal1 217 259 217 259 1 vdd
rlabel metal1 251 200 251 200 1 c4
rlabel metal1 82 200 82 200 1 g3_bar
rlabel metal1 80 194 80 194 1 vdd
rlabel metal1 88 108 88 108 1 gnd
rlabel metal1 62 128 62 128 1 p4_bar
rlabel metal1 89 102 89 102 1 vdd
rlabel metal1 94 18 94 18 1 gnd
rlabel metal1 52 9 52 9 1 g4_bar
rlabel metal1 173 160 173 160 1 vdd
rlabel metal1 175 88 175 88 1 gnd
rlabel metal1 133 9 133 9 1 gnd
rlabel metal1 144 81 144 81 1 vdd
rlabel metal1 236 23 236 23 1 gnd
rlabel metal1 232 107 232 107 1 vdd
rlabel metal1 266 48 266 48 7 c5
rlabel metal1 33 706 33 706 5 vdd
rlabel metal1 34 624 34 624 1 gnd
rlabel metal1 15 617 15 617 1 b1
rlabel metal1 9 617 9 617 3 a1
rlabel metal1 71 763 71 763 5 vdd
rlabel metal1 61 691 61 691 1 gnd
rlabel metal1 55 725 55 725 1 a0
rlabel metal1 55 718 55 718 1 b0
rlabel metal1 52 391 52 391 1 g2_bar
rlabel metal1 28 532 28 532 1 vdd
rlabel metal1 29 449 29 449 1 gnd
rlabel metal1 10 441 10 441 1 b2
rlabel metal1 4 441 4 441 3 a2
rlabel metal1 57 319 57 319 1 p3_bar
rlabel metal1 26 359 26 359 1 vdd
rlabel metal1 28 276 28 276 1 gnd
rlabel metal1 10 274 10 274 1 b3
rlabel metal1 3 274 3 274 3 a3
rlabel metal1 26 158 26 158 1 vdd
rlabel metal1 30 76 30 76 1 gnd
rlabel metal1 11 72 11 72 1 b4
rlabel metal1 5 72 5 72 3 a4
rlabel metal1 239 706 239 706 1 gnd
rlabel metal1 223 855 223 855 5 vdd
rlabel metal1 273 732 273 732 1 s0
rlabel metal1 326 746 326 746 1 vdd
rlabel metal1 337 597 337 597 1 gnd
rlabel metal1 374 624 374 624 7 p1
rlabel metal1 449 630 449 630 7 s1
rlabel metal1 417 603 417 603 1 gnd
rlabel metal1 406 753 406 753 1 vdd
rlabel metal1 324 575 324 575 1 vdd
rlabel metal1 339 425 339 425 1 gnd
rlabel metal1 369 452 369 452 1 p2
rlabel metal1 430 425 430 425 1 gnd
rlabel metal1 418 575 418 575 1 vdd
rlabel metal1 332 408 332 408 1 vdd
rlabel metal1 327 259 327 259 1 gnd
rlabel metal1 374 286 374 286 1 p3
rlabel metal1 416 260 416 260 1 gnd
rlabel metal1 417 408 417 408 1 vdd
rlabel metal1 460 287 460 287 7 s3
rlabel metal1 335 204 335 204 1 vdd
rlabel metal1 343 54 343 54 1 gnd
rlabel metal1 375 81 375 81 1 p4
rlabel metal1 414 245 414 245 1 vdd
rlabel metal1 428 96 428 96 1 gnd
rlabel metal1 456 123 456 123 1 s4
rlabel metal1 459 452 459 452 7 s2
rlabel metal1 207 765 207 765 1 vdd
rlabel metal1 310 657 310 657 1 vdd
rlabel metal1 389 663 389 663 1 vdd
rlabel metal1 309 484 309 484 1 vdd
rlabel metal1 399 484 399 484 1 vdd
rlabel metal1 313 319 313 319 1 vdd
rlabel metal1 400 319 400 319 1 vdd
rlabel metal1 314 114 314 114 1 vdd
rlabel metal1 397 155 397 155 1 vdd
rlabel metal2 327 852 327 852 1 clk
rlabel metal1 338 860 338 860 5 vdd
rlabel metal1 356 758 356 758 1 gnd
rlabel metal1 416 810 416 810 1 S0_out
rlabel metal2 -76 865 -76 865 1 clk
rlabel metal1 -69 873 -69 873 5 vdd
rlabel metal1 -57 771 -57 771 1 gnd
rlabel metal1 -52 660 -52 660 1 gnd
rlabel metal2 -76 755 -76 755 1 clk
rlabel metal1 -58 763 -58 763 1 vdd
rlabel metal1 -104 697 -104 697 3 B0_in
rlabel metal2 -189 695 -189 695 1 clk
rlabel metal1 -175 703 -175 703 1 vdd
rlabel metal1 -173 600 -173 600 1 gnd
rlabel metal1 -216 637 -216 637 3 B1_in
rlabel metal1 -66 521 -66 521 1 gnd
rlabel metal2 -85 615 -85 615 1 clk
rlabel metal1 -72 624 -72 624 1 vdd
rlabel metal1 -116 558 -116 558 1 A1_in
rlabel metal1 -185 562 -185 562 1 vdd
rlabel metal2 -197 553 -197 553 1 clk
rlabel metal1 -183 459 -183 459 1 gnd
rlabel metal1 -225 495 -225 495 3 B2_in
rlabel metal1 -61 462 -61 462 1 vdd
rlabel metal2 -88 454 -88 454 1 clk
rlabel metal1 -71 360 -71 360 1 gnd
rlabel metal1 -121 396 -121 396 1 A2_in
rlabel metal1 -192 408 -192 408 1 vdd
rlabel metal1 -195 306 -195 306 1 gnd
rlabel metal2 -212 400 -212 400 1 clk
rlabel metal1 -241 342 -241 342 3 B3_in
rlabel metal1 -75 289 -75 289 1 vdd
rlabel metal2 -95 282 -95 282 1 clk
rlabel metal1 -75 188 -75 188 1 gnd
rlabel metal1 -128 223 -128 223 1 A3_in
rlabel metal1 -200 178 -200 178 1 vdd
rlabel metal1 -198 76 -198 76 1 gnd
rlabel metal2 -213 170 -213 170 1 clk
rlabel metal1 -247 112 -247 112 3 B4_in
rlabel metal1 -74 -11 -74 -11 1 gnd
rlabel metal1 -77 91 -77 91 1 vdd
rlabel metal1 -134 25 -134 25 1 A4_in
rlabel metal1 507 706 507 706 1 vdd
rlabel metal2 484 697 484 697 1 clk
rlabel metal1 504 604 504 604 1 gnd
rlabel metal1 571 656 571 656 7 S1_out
rlabel metal1 512 528 512 528 1 vdd
rlabel metal1 515 425 515 425 1 gnd
rlabel metal2 497 519 497 519 1 clk
rlabel metal1 506 370 506 370 1 vdd
rlabel metal2 497 362 497 362 1 clk
rlabel metal1 504 268 504 268 1 gnd
rlabel metal1 582 478 582 478 7 S2_out
rlabel metal1 585 320 585 320 7 S3_out
rlabel metal1 513 149 513 149 1 gnd
rlabel metal1 515 252 515 252 1 vdd
rlabel metal2 497 243 497 243 1 clk
rlabel metal1 583 202 583 202 1 S4_out
rlabel metal1 520 129 520 129 1 vdd
rlabel metal1 516 26 516 26 1 gnd
rlabel metal2 500 120 500 120 1 clk
rlabel metal1 589 79 589 79 7 COUT_out
rlabel metal2 -98 83 -98 83 1 clk
rlabel metal1 -104 808 -104 808 1 A0_in
<< end >>
