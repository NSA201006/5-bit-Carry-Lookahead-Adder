magic
tech scmos
timestamp 1762626811
<< nwell >>
rect -12 2 53 34
rect -12 -18 18 2
rect 72 -2 98 30
<< ntransistor >>
rect -1 -34 1 -24
rect 31 -48 33 -8
rect 37 -48 39 -8
rect 55 -28 57 -8
rect 64 -28 66 -8
rect 83 -20 85 -10
<< ptransistor >>
rect -1 -12 1 28
rect 5 -12 7 28
rect 21 8 23 28
rect 37 8 39 28
rect 83 4 85 24
<< ndiffusion >>
rect 30 -12 31 -8
rect -6 -30 -1 -24
rect -2 -34 -1 -30
rect 1 -28 2 -24
rect 1 -34 6 -28
rect 26 -48 31 -12
rect 33 -48 37 -8
rect 39 -44 44 -8
rect 52 -12 55 -8
rect 48 -28 55 -12
rect 57 -28 64 -8
rect 66 -24 74 -8
rect 78 -16 83 -10
rect 82 -20 83 -16
rect 85 -14 88 -10
rect 85 -20 92 -14
rect 66 -28 70 -24
rect 39 -48 40 -44
<< pdiffusion >>
rect -2 24 -1 28
rect -6 -12 -1 24
rect 1 -12 5 28
rect 7 -8 12 28
rect 20 24 21 28
rect 16 8 21 24
rect 23 12 28 28
rect 23 8 24 12
rect 36 24 37 28
rect 32 8 37 24
rect 39 12 44 28
rect 39 8 40 12
rect 82 20 83 24
rect 78 4 83 20
rect 85 8 92 24
rect 85 4 88 8
rect 7 -12 8 -8
<< ndcontact >>
rect 26 -12 30 -8
rect -6 -34 -2 -30
rect 2 -28 6 -24
rect 48 -12 52 -8
rect 78 -20 82 -16
rect 88 -14 92 -10
rect 70 -28 74 -24
rect 40 -48 44 -44
<< pdcontact >>
rect -6 24 -2 28
rect 16 24 20 28
rect 24 8 28 12
rect 32 24 36 28
rect 40 8 44 12
rect 78 20 82 24
rect 88 4 92 8
rect 8 -12 12 -8
<< polysilicon >>
rect -1 28 1 31
rect 5 28 7 35
rect 21 28 23 40
rect 37 28 39 31
rect 83 24 85 32
rect 21 5 23 8
rect 37 3 39 8
rect 31 -8 33 -5
rect 83 -3 85 4
rect 37 -8 39 -7
rect 55 -8 57 -7
rect 64 -8 66 -5
rect -1 -24 1 -12
rect 5 -15 7 -12
rect -1 -37 1 -34
rect 83 -10 85 -7
rect 83 -23 85 -20
rect 55 -31 57 -28
rect 64 -31 66 -28
rect 31 -49 33 -48
rect 37 -51 39 -48
<< polycontact >>
rect 33 3 37 7
rect 81 -7 85 -3
rect -5 -23 -1 -19
rect 64 -35 68 -31
rect 29 -53 33 -49
<< metal1 >>
rect -6 43 81 46
rect -6 28 -2 43
rect 16 28 20 43
rect 32 28 36 43
rect 78 24 81 43
rect 44 11 53 12
rect 44 8 77 11
rect 24 7 28 8
rect 24 3 33 7
rect 24 0 28 3
rect 20 -3 30 0
rect -9 -23 -5 -19
rect 8 -21 12 -12
rect 2 -24 12 -21
rect -6 -56 -2 -34
rect 9 -50 12 -24
rect 20 -31 23 -3
rect 26 -8 30 -3
rect 48 -8 51 8
rect 74 -3 77 8
rect 88 -3 92 4
rect 74 -6 81 -3
rect 88 -7 94 -3
rect 88 -10 92 -7
rect 20 -35 64 -31
rect 9 -53 29 -50
rect 40 -56 44 -48
rect 71 -56 74 -28
rect 78 -56 81 -20
rect -6 -59 81 -56
<< pm12contact >>
rect 5 35 10 40
rect 23 35 28 40
rect 37 -7 42 -2
rect 55 -7 60 -2
<< metal2 >>
rect 10 35 23 38
rect 13 -4 16 35
rect 13 -7 37 -4
rect 42 -7 55 -4
<< labels >>
rlabel metal1 -7 -21 -7 -21 3 D
rlabel metal1 9 45 9 45 5 vdd
rlabel metal2 12 36 12 36 1 clk
rlabel metal1 10 -20 10 -20 1 X
rlabel metal1 54 10 54 10 7 Q_bar
rlabel metal1 28 -3 28 -3 1 Y
rlabel metal1 20 -58 20 -58 1 gnd
rlabel metal1 93 -5 93 -5 7 Q
<< end >>
