magic
tech scmos
timestamp 1764616678
<< nwell >>
rect -1 53 23 85
rect -11 -37 13 -5
rect 29 -31 53 1
<< ntransistor >>
rect 10 37 12 47
rect -4 5 -2 25
rect 25 8 27 28
rect 0 -53 2 -43
rect 40 -57 42 -37
<< ptransistor >>
rect 10 59 12 79
rect 0 -31 2 -11
rect 40 -25 42 -5
<< ndiffusion >>
rect 5 41 10 47
rect 9 37 10 41
rect 12 43 13 47
rect 12 37 17 43
rect -10 10 -4 25
rect -5 5 -4 10
rect -2 9 3 25
rect -2 5 -1 9
rect 19 13 25 28
rect 24 8 25 13
rect 27 12 32 28
rect 27 8 28 12
rect -5 -49 0 -43
rect -1 -53 0 -49
rect 2 -47 3 -43
rect 2 -53 7 -47
rect 35 -53 40 -37
rect 39 -57 40 -53
rect 42 -41 43 -37
rect 42 -57 47 -41
<< pdiffusion >>
rect 9 75 10 79
rect 5 59 10 75
rect 12 63 17 79
rect 12 59 13 63
rect 39 -9 40 -5
rect -1 -15 0 -11
rect -5 -31 0 -15
rect 2 -27 7 -11
rect 35 -25 40 -9
rect 42 -21 47 -5
rect 42 -25 43 -21
rect 2 -31 3 -27
<< ndcontact >>
rect 5 37 9 41
rect 13 43 17 47
rect -1 5 3 9
rect 28 8 32 12
rect -5 -53 -1 -49
rect 3 -47 7 -43
rect 35 -57 39 -53
rect 43 -41 47 -37
<< pdcontact >>
rect 5 75 9 79
rect 13 59 17 63
rect 35 -9 39 -5
rect -5 -15 -1 -11
rect 43 -25 47 -21
rect 3 -31 7 -27
<< polysilicon >>
rect 10 79 12 82
rect 10 47 12 59
rect 10 34 12 37
rect 25 28 27 29
rect -4 25 -2 26
rect 25 5 27 8
rect -4 2 -2 5
rect 40 -5 42 -2
rect 0 -11 2 -8
rect 0 -43 2 -31
rect 40 -37 42 -25
rect 0 -56 2 -53
rect 40 -60 42 -57
<< polycontact >>
rect 6 48 10 52
rect -6 26 -2 30
rect 23 29 27 33
rect -4 -42 0 -38
<< polynpluscontact >>
rect 36 -36 40 -32
<< metal1 >>
rect -16 86 38 89
rect -16 -1 -13 86
rect 5 79 8 86
rect -10 48 6 51
rect 14 51 17 59
rect 14 48 26 51
rect -10 30 -7 48
rect 14 47 17 48
rect 5 33 8 37
rect 23 33 26 48
rect 5 30 10 33
rect -10 27 -6 30
rect 29 5 32 8
rect 0 2 32 5
rect -16 -4 0 -1
rect -5 -11 -2 -4
rect -11 -42 -4 -39
rect 4 -39 7 -31
rect 29 -33 32 2
rect 35 -5 38 86
rect 29 -36 36 -33
rect 44 -33 47 -25
rect 44 -36 53 -33
rect 44 -37 47 -36
rect 4 -42 19 -39
rect 4 -43 7 -42
rect -5 -60 -2 -53
rect 35 -60 38 -57
rect -5 -63 10 -60
rect 15 -63 38 -60
<< m2contact >>
rect 10 28 15 33
rect -16 -44 -11 -39
rect 19 -42 24 -37
rect 10 -65 15 -60
<< ndm12contact >>
rect -10 5 -5 10
rect 19 8 24 13
<< metal2 >>
rect -16 5 -10 10
rect -16 -39 -13 5
rect 12 -60 15 28
rect 19 -37 22 8
<< labels >>
rlabel metal1 10 -40 10 -40 1 A_bar
rlabel metal1 4 88 4 88 4 vdd
rlabel metal1 -5 49 -5 49 1 B
rlabel metal1 20 49 20 49 7 B_bar
rlabel metal1 31 3 31 3 7 Y_bar
rlabel metal1 50 -35 50 -35 7 Y
rlabel metal1 1 -62 1 -62 1 gnd
rlabel metal1 -10 -41 -10 -41 1 A
<< end >>
