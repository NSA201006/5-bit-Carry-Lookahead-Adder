magic
tech scmos
timestamp 1764345749
<< nwell >>
rect 172 848 237 880
rect 172 828 202 848
rect 256 844 282 876
rect 489 837 513 869
rect 575 835 640 867
rect 575 815 605 835
rect 659 831 685 863
rect 172 737 237 769
rect 172 717 202 737
rect 256 733 282 765
rect 327 746 361 778
rect 479 747 503 779
rect 519 753 543 785
rect 59 677 124 709
rect 59 657 89 677
rect 143 673 169 705
rect 290 669 324 721
rect 368 714 392 746
rect 592 729 616 761
rect 671 735 695 767
rect 358 664 394 684
rect 358 632 418 664
rect 582 639 606 671
rect 622 645 646 677
rect 661 645 685 677
rect 701 651 725 683
rect 733 680 798 712
rect 733 660 763 680
rect 817 676 843 708
rect 162 598 227 630
rect 162 578 192 598
rect 246 594 272 626
rect 425 607 459 639
rect 290 569 324 601
rect 51 536 116 568
rect 51 516 81 536
rect 135 532 161 564
rect 285 495 319 547
rect 358 534 394 586
rect 590 557 614 589
rect 681 557 705 589
rect 417 522 475 554
rect 348 476 384 496
rect 160 437 225 469
rect 160 417 190 437
rect 244 433 270 465
rect 348 444 408 476
rect 471 471 507 491
rect 36 383 101 415
rect 36 363 66 383
rect 120 379 146 411
rect 285 395 319 427
rect 422 420 456 452
rect 471 439 531 471
rect 580 467 604 499
rect 620 473 644 505
rect 671 467 695 499
rect 711 473 735 505
rect 745 502 810 534
rect 745 482 775 502
rect 829 498 855 530
rect 284 322 318 374
rect 339 346 375 398
rect 595 391 619 423
rect 682 391 706 423
rect 461 327 519 359
rect 745 345 810 377
rect 153 264 218 296
rect 153 244 183 264
rect 237 260 263 292
rect 346 285 382 305
rect 585 301 609 333
rect 625 307 649 339
rect 672 301 696 333
rect 712 307 736 339
rect 745 325 775 345
rect 829 341 855 373
rect 284 222 318 254
rect 346 253 406 285
rect 422 228 456 260
rect 466 254 502 274
rect 466 222 526 254
rect 679 228 703 260
rect 745 226 810 258
rect 35 153 100 185
rect 35 133 65 153
rect 119 149 145 181
rect 286 122 320 174
rect 346 155 382 207
rect 597 186 621 218
rect 745 206 775 226
rect 829 222 855 254
rect 424 143 482 175
rect 669 138 693 170
rect 709 144 733 176
rect 150 66 215 98
rect 340 97 376 117
rect 482 102 518 122
rect 340 96 400 97
rect 150 46 180 66
rect 234 62 260 94
rect 340 65 434 96
rect 482 70 542 102
rect 587 96 611 128
rect 627 102 651 134
rect 748 103 813 135
rect 748 83 778 103
rect 832 99 858 131
rect 400 64 434 65
rect 286 22 320 54
<< ntransistor >>
rect 183 812 185 822
rect 215 798 217 838
rect 221 798 223 838
rect 239 818 241 838
rect 248 818 250 838
rect 267 826 269 836
rect 500 821 502 831
rect 486 789 488 809
rect 515 792 517 812
rect 586 799 588 809
rect 618 785 620 825
rect 624 785 626 825
rect 642 805 644 825
rect 651 805 653 825
rect 670 813 672 823
rect 183 701 185 711
rect 215 687 217 727
rect 221 687 223 727
rect 239 707 241 727
rect 248 707 250 727
rect 267 715 269 725
rect 338 713 340 733
rect 348 713 350 733
rect 490 731 492 741
rect 530 727 532 747
rect 603 713 605 723
rect 682 719 684 729
rect 379 698 381 708
rect 589 681 591 701
rect 618 684 620 704
rect 668 687 670 707
rect 697 690 699 710
rect 70 641 72 651
rect 102 627 104 667
rect 108 627 110 667
rect 126 647 128 667
rect 135 647 137 667
rect 154 655 156 665
rect 301 646 303 656
rect 311 646 313 656
rect 301 615 303 635
rect 311 615 313 635
rect 370 610 372 620
rect 380 610 382 620
rect 405 614 407 624
rect 593 623 595 633
rect 633 619 635 639
rect 672 629 674 639
rect 712 625 714 645
rect 744 644 746 654
rect 776 630 778 670
rect 782 630 784 670
rect 800 650 802 670
rect 809 650 811 670
rect 828 658 830 668
rect 173 562 175 572
rect 205 548 207 588
rect 211 548 213 588
rect 229 568 231 588
rect 238 568 240 588
rect 257 576 259 586
rect 62 500 64 510
rect 94 486 96 526
rect 100 486 102 526
rect 118 506 120 526
rect 127 506 129 526
rect 146 514 148 524
rect 436 574 438 594
rect 446 574 448 594
rect 601 541 603 551
rect 692 541 694 551
rect 370 512 372 522
rect 380 512 382 522
rect 296 472 298 482
rect 306 472 308 482
rect 296 441 298 461
rect 306 441 308 461
rect 428 489 430 509
rect 438 489 440 509
rect 462 506 464 516
rect 587 509 589 529
rect 616 512 618 532
rect 678 509 680 529
rect 707 512 709 532
rect 171 401 173 411
rect 203 387 205 427
rect 209 387 211 427
rect 227 407 229 427
rect 236 407 238 427
rect 255 415 257 425
rect 360 422 362 432
rect 370 422 372 432
rect 395 426 397 436
rect 591 451 593 461
rect 631 447 633 467
rect 682 451 684 461
rect 722 447 724 467
rect 756 466 758 476
rect 788 452 790 492
rect 794 452 796 492
rect 812 472 814 492
rect 821 472 823 492
rect 840 480 842 490
rect 483 417 485 427
rect 493 417 495 427
rect 518 421 520 431
rect 47 347 49 357
rect 79 333 81 373
rect 85 333 87 373
rect 103 353 105 373
rect 112 353 114 373
rect 131 361 133 371
rect 433 387 435 407
rect 443 387 445 407
rect 606 375 608 385
rect 693 375 695 385
rect 351 324 353 334
rect 361 324 363 334
rect 592 343 594 363
rect 621 346 623 366
rect 679 343 681 363
rect 708 346 710 366
rect 295 299 297 309
rect 305 299 307 309
rect 295 268 297 288
rect 305 268 307 288
rect 164 228 166 238
rect 196 214 198 254
rect 202 214 204 254
rect 220 234 222 254
rect 229 234 231 254
rect 248 242 250 252
rect 472 294 474 314
rect 482 294 484 314
rect 506 311 508 321
rect 596 285 598 295
rect 636 281 638 301
rect 756 309 758 319
rect 683 285 685 295
rect 723 281 725 301
rect 788 295 790 335
rect 794 295 796 335
rect 812 315 814 335
rect 821 315 823 335
rect 840 323 842 333
rect 358 231 360 241
rect 368 231 370 241
rect 393 235 395 245
rect 46 117 48 127
rect 78 103 80 143
rect 84 103 86 143
rect 102 123 104 143
rect 111 123 113 143
rect 130 131 132 141
rect 433 195 435 215
rect 443 195 445 215
rect 478 200 480 210
rect 488 200 490 210
rect 513 204 515 214
rect 690 212 692 222
rect 676 180 678 200
rect 705 183 707 203
rect 756 190 758 200
rect 608 170 610 180
rect 788 176 790 216
rect 794 176 796 216
rect 812 196 814 216
rect 821 196 823 216
rect 840 204 842 214
rect 358 133 360 143
rect 368 133 370 143
rect 594 138 596 158
rect 623 141 625 161
rect 297 99 299 109
rect 307 99 309 109
rect 297 68 299 88
rect 307 68 309 88
rect 435 110 437 130
rect 445 110 447 130
rect 469 127 471 137
rect 161 30 163 40
rect 193 16 195 56
rect 199 16 201 56
rect 217 36 219 56
rect 226 36 228 56
rect 245 44 247 54
rect 680 122 682 132
rect 720 118 722 138
rect 598 80 600 90
rect 638 76 640 96
rect 352 43 354 53
rect 362 43 364 53
rect 387 47 389 57
rect 759 67 761 77
rect 411 31 413 51
rect 421 31 423 51
rect 494 48 496 58
rect 504 48 506 58
rect 529 52 531 62
rect 791 53 793 93
rect 797 53 799 93
rect 815 73 817 93
rect 824 73 826 93
rect 843 81 845 91
<< ptransistor >>
rect 183 834 185 874
rect 189 834 191 874
rect 205 854 207 874
rect 221 854 223 874
rect 267 850 269 870
rect 500 843 502 863
rect 586 821 588 861
rect 592 821 594 861
rect 608 841 610 861
rect 624 841 626 861
rect 670 837 672 857
rect 183 723 185 763
rect 189 723 191 763
rect 205 743 207 763
rect 221 743 223 763
rect 267 739 269 759
rect 338 752 340 772
rect 348 752 350 772
rect 490 753 492 773
rect 530 759 532 779
rect 70 663 72 703
rect 76 663 78 703
rect 92 683 94 703
rect 108 683 110 703
rect 154 679 156 699
rect 301 675 303 715
rect 311 675 313 715
rect 379 720 381 740
rect 603 735 605 755
rect 682 741 684 761
rect 370 638 372 678
rect 380 638 382 678
rect 405 638 407 658
rect 593 645 595 665
rect 633 651 635 671
rect 672 651 674 671
rect 712 657 714 677
rect 744 666 746 706
rect 750 666 752 706
rect 766 686 768 706
rect 782 686 784 706
rect 828 682 830 702
rect 173 584 175 624
rect 179 584 181 624
rect 195 604 197 624
rect 211 604 213 624
rect 257 600 259 620
rect 436 613 438 633
rect 446 613 448 633
rect 62 522 64 562
rect 68 522 70 562
rect 84 542 86 562
rect 100 542 102 562
rect 146 538 148 558
rect 301 575 303 595
rect 311 575 313 595
rect 296 501 298 541
rect 306 501 308 541
rect 370 540 372 580
rect 380 540 382 580
rect 601 563 603 583
rect 692 563 694 583
rect 428 528 430 548
rect 438 528 440 548
rect 462 528 464 548
rect 171 423 173 463
rect 177 423 179 463
rect 193 443 195 463
rect 209 443 211 463
rect 255 439 257 459
rect 360 450 362 490
rect 370 450 372 490
rect 395 450 397 470
rect 47 369 49 409
rect 53 369 55 409
rect 69 389 71 409
rect 85 389 87 409
rect 131 385 133 405
rect 433 426 435 446
rect 443 426 445 446
rect 483 445 485 485
rect 493 445 495 485
rect 591 473 593 493
rect 631 479 633 499
rect 518 445 520 465
rect 682 473 684 493
rect 722 479 724 499
rect 756 488 758 528
rect 762 488 764 528
rect 778 508 780 528
rect 794 508 796 528
rect 840 504 842 524
rect 296 401 298 421
rect 306 401 308 421
rect 295 328 297 368
rect 305 328 307 368
rect 351 352 353 392
rect 361 352 363 392
rect 606 397 608 417
rect 693 397 695 417
rect 472 333 474 353
rect 482 333 484 353
rect 506 333 508 353
rect 164 250 166 290
rect 170 250 172 290
rect 186 270 188 290
rect 202 270 204 290
rect 248 266 250 286
rect 358 259 360 299
rect 368 259 370 299
rect 596 307 598 327
rect 636 313 638 333
rect 683 307 685 327
rect 723 313 725 333
rect 756 331 758 371
rect 762 331 764 371
rect 778 351 780 371
rect 794 351 796 371
rect 840 347 842 367
rect 393 259 395 279
rect 295 228 297 248
rect 305 228 307 248
rect 433 234 435 254
rect 443 234 445 254
rect 478 228 480 268
rect 488 228 490 268
rect 513 228 515 248
rect 690 234 692 254
rect 46 139 48 179
rect 52 139 54 179
rect 68 159 70 179
rect 84 159 86 179
rect 130 155 132 175
rect 297 128 299 168
rect 307 128 309 168
rect 358 161 360 201
rect 368 161 370 201
rect 756 212 758 252
rect 762 212 764 252
rect 778 232 780 252
rect 794 232 796 252
rect 840 228 842 248
rect 608 192 610 212
rect 435 149 437 169
rect 445 149 447 169
rect 469 149 471 169
rect 680 144 682 164
rect 720 150 722 170
rect 161 52 163 92
rect 167 52 169 92
rect 183 72 185 92
rect 199 72 201 92
rect 245 68 247 88
rect 352 71 354 111
rect 362 71 364 111
rect 387 71 389 91
rect 411 70 413 90
rect 421 70 423 90
rect 494 76 496 116
rect 504 76 506 116
rect 598 102 600 122
rect 638 108 640 128
rect 529 76 531 96
rect 759 89 761 129
rect 765 89 767 129
rect 781 109 783 129
rect 797 109 799 129
rect 843 105 845 125
rect 297 28 299 48
rect 307 28 309 48
<< ndiffusion >>
rect 214 834 215 838
rect 178 816 183 822
rect 182 812 183 816
rect 185 818 186 822
rect 185 812 190 818
rect 210 798 215 834
rect 217 798 221 838
rect 223 802 228 838
rect 236 834 239 838
rect 232 818 239 834
rect 241 818 248 838
rect 250 822 258 838
rect 262 830 267 836
rect 266 826 267 830
rect 269 832 272 836
rect 269 826 276 832
rect 495 825 500 831
rect 250 818 254 822
rect 499 821 500 825
rect 502 827 503 831
rect 502 821 507 827
rect 617 821 618 825
rect 223 798 224 802
rect 480 794 486 809
rect 485 789 486 794
rect 488 793 493 809
rect 488 789 489 793
rect 509 797 515 812
rect 514 792 515 797
rect 517 796 522 812
rect 581 803 586 809
rect 585 799 586 803
rect 588 805 589 809
rect 588 799 593 805
rect 517 792 518 796
rect 613 785 618 821
rect 620 785 624 825
rect 626 789 631 825
rect 639 821 642 825
rect 635 805 642 821
rect 644 805 651 825
rect 653 809 661 825
rect 665 817 670 823
rect 669 813 670 817
rect 672 819 675 823
rect 672 813 679 819
rect 653 805 657 809
rect 626 785 627 789
rect 214 723 215 727
rect 178 705 183 711
rect 182 701 183 705
rect 185 707 186 711
rect 185 701 190 707
rect 210 687 215 723
rect 217 687 221 727
rect 223 691 228 727
rect 236 723 239 727
rect 232 707 239 723
rect 241 707 248 727
rect 250 711 258 727
rect 262 719 267 725
rect 266 715 267 719
rect 269 721 272 725
rect 269 715 276 721
rect 333 717 338 733
rect 250 707 254 711
rect 223 687 224 691
rect 337 713 338 717
rect 340 713 348 733
rect 350 729 351 733
rect 350 713 355 729
rect 485 735 490 741
rect 489 731 490 735
rect 492 737 493 741
rect 492 731 497 737
rect 525 731 530 747
rect 529 727 530 731
rect 532 743 533 747
rect 532 727 537 743
rect 677 723 682 729
rect 598 717 603 723
rect 602 713 603 717
rect 605 719 606 723
rect 681 719 682 723
rect 684 725 685 729
rect 684 719 689 725
rect 605 713 610 719
rect 374 702 379 708
rect 378 698 379 702
rect 381 704 382 708
rect 381 698 386 704
rect 583 686 589 701
rect 588 681 589 686
rect 591 685 596 701
rect 591 681 592 685
rect 612 689 618 704
rect 617 684 618 689
rect 620 688 625 704
rect 620 684 621 688
rect 662 692 668 707
rect 667 687 668 692
rect 670 691 675 707
rect 670 687 671 691
rect 691 695 697 710
rect 696 690 697 695
rect 699 694 704 710
rect 699 690 700 694
rect 101 663 102 667
rect 65 645 70 651
rect 69 641 70 645
rect 72 647 73 651
rect 72 641 77 647
rect 97 627 102 663
rect 104 627 108 667
rect 110 631 115 667
rect 123 663 126 667
rect 119 647 126 663
rect 128 647 135 667
rect 137 651 145 667
rect 149 659 154 665
rect 153 655 154 659
rect 156 661 159 665
rect 156 655 163 661
rect 137 647 141 651
rect 296 650 301 656
rect 300 646 301 650
rect 303 652 305 656
rect 309 652 311 656
rect 303 646 311 652
rect 313 650 318 656
rect 313 646 314 650
rect 775 666 776 670
rect 110 627 111 631
rect 300 631 301 635
rect 296 615 301 631
rect 303 615 311 635
rect 313 619 318 635
rect 739 648 744 654
rect 313 615 314 619
rect 365 614 370 620
rect 369 610 370 614
rect 372 616 374 620
rect 378 616 380 620
rect 372 610 380 616
rect 382 614 387 620
rect 400 618 405 624
rect 404 614 405 618
rect 407 620 408 624
rect 407 614 412 620
rect 382 610 383 614
rect 588 627 593 633
rect 592 623 593 627
rect 595 629 596 633
rect 595 623 600 629
rect 628 623 633 639
rect 632 619 633 623
rect 635 635 636 639
rect 635 619 640 635
rect 667 633 672 639
rect 671 629 672 633
rect 674 635 675 639
rect 674 629 679 635
rect 707 629 712 645
rect 711 625 712 629
rect 714 641 715 645
rect 743 644 744 648
rect 746 650 747 654
rect 746 644 751 650
rect 714 625 719 641
rect 771 630 776 666
rect 778 630 782 670
rect 784 634 789 670
rect 797 666 800 670
rect 793 650 800 666
rect 802 650 809 670
rect 811 654 819 670
rect 823 662 828 668
rect 827 658 828 662
rect 830 664 833 668
rect 830 658 837 664
rect 811 650 815 654
rect 784 630 785 634
rect 204 584 205 588
rect 168 566 173 572
rect 172 562 173 566
rect 175 568 176 572
rect 175 562 180 568
rect 200 548 205 584
rect 207 548 211 588
rect 213 552 218 588
rect 226 584 229 588
rect 222 568 229 584
rect 231 568 238 588
rect 240 572 248 588
rect 252 580 257 586
rect 256 576 257 580
rect 259 582 262 586
rect 259 576 266 582
rect 240 568 244 572
rect 213 548 214 552
rect 93 522 94 526
rect 57 504 62 510
rect 61 500 62 504
rect 64 506 65 510
rect 64 500 69 506
rect 89 486 94 522
rect 96 486 100 526
rect 102 490 107 526
rect 115 522 118 526
rect 111 506 118 522
rect 120 506 127 526
rect 129 510 137 526
rect 141 518 146 524
rect 145 514 146 518
rect 148 520 151 524
rect 148 514 155 520
rect 129 506 133 510
rect 431 578 436 594
rect 435 574 436 578
rect 438 574 446 594
rect 448 590 449 594
rect 448 574 453 590
rect 596 545 601 551
rect 600 541 601 545
rect 603 547 604 551
rect 603 541 608 547
rect 687 545 692 551
rect 691 541 692 545
rect 694 547 695 551
rect 694 541 699 547
rect 365 516 370 522
rect 369 512 370 516
rect 372 518 374 522
rect 378 518 380 522
rect 372 512 380 518
rect 382 516 387 522
rect 382 512 383 516
rect 457 510 462 516
rect 102 486 103 490
rect 423 493 428 509
rect 291 476 296 482
rect 295 472 296 476
rect 298 478 300 482
rect 304 478 306 482
rect 298 472 306 478
rect 308 476 313 482
rect 308 472 309 476
rect 295 457 296 461
rect 291 441 296 457
rect 298 441 306 461
rect 308 445 313 461
rect 427 489 428 493
rect 430 489 438 509
rect 440 505 441 509
rect 461 506 462 510
rect 464 512 465 516
rect 464 506 469 512
rect 581 514 587 529
rect 586 509 587 514
rect 589 513 594 529
rect 589 509 590 513
rect 610 517 616 532
rect 615 512 616 517
rect 618 516 623 532
rect 618 512 619 516
rect 672 514 678 529
rect 677 509 678 514
rect 680 513 685 529
rect 680 509 681 513
rect 701 517 707 532
rect 706 512 707 517
rect 709 516 714 532
rect 709 512 710 516
rect 440 489 445 505
rect 308 441 309 445
rect 202 423 203 427
rect 166 405 171 411
rect 170 401 171 405
rect 173 407 174 411
rect 173 401 178 407
rect 198 387 203 423
rect 205 387 209 427
rect 211 391 216 427
rect 224 423 227 427
rect 220 407 227 423
rect 229 407 236 427
rect 238 411 246 427
rect 250 419 255 425
rect 254 415 255 419
rect 257 421 260 425
rect 355 426 360 432
rect 359 422 360 426
rect 362 428 364 432
rect 368 428 370 432
rect 362 422 370 428
rect 372 426 377 432
rect 390 430 395 436
rect 394 426 395 430
rect 397 432 398 436
rect 397 426 402 432
rect 787 488 788 492
rect 586 455 591 461
rect 590 451 591 455
rect 593 457 594 461
rect 593 451 598 457
rect 626 451 631 467
rect 630 447 631 451
rect 633 463 634 467
rect 633 447 638 463
rect 751 470 756 476
rect 677 455 682 461
rect 681 451 682 455
rect 684 457 685 461
rect 684 451 689 457
rect 717 451 722 467
rect 721 447 722 451
rect 724 463 725 467
rect 755 466 756 470
rect 758 472 759 476
rect 758 466 763 472
rect 724 447 729 463
rect 783 452 788 488
rect 790 452 794 492
rect 796 456 801 492
rect 809 488 812 492
rect 805 472 812 488
rect 814 472 821 492
rect 823 476 831 492
rect 835 484 840 490
rect 839 480 840 484
rect 842 486 845 490
rect 842 480 849 486
rect 823 472 827 476
rect 796 452 797 456
rect 372 422 373 426
rect 257 415 264 421
rect 238 407 242 411
rect 478 421 483 427
rect 482 417 483 421
rect 485 423 487 427
rect 491 423 493 427
rect 485 417 493 423
rect 495 421 500 427
rect 513 425 518 431
rect 517 421 518 425
rect 520 427 521 431
rect 520 421 525 427
rect 495 417 496 421
rect 211 387 212 391
rect 78 369 79 373
rect 42 351 47 357
rect 46 347 47 351
rect 49 353 50 357
rect 49 347 54 353
rect 74 333 79 369
rect 81 333 85 373
rect 87 337 92 373
rect 100 369 103 373
rect 96 353 103 369
rect 105 353 112 373
rect 114 357 122 373
rect 126 365 131 371
rect 130 361 131 365
rect 133 367 136 371
rect 133 361 140 367
rect 114 353 118 357
rect 87 333 88 337
rect 428 391 433 407
rect 432 387 433 391
rect 435 387 443 407
rect 445 403 446 407
rect 445 387 450 403
rect 601 379 606 385
rect 605 375 606 379
rect 608 381 609 385
rect 608 375 613 381
rect 688 379 693 385
rect 692 375 693 379
rect 695 381 696 385
rect 695 375 700 381
rect 346 328 351 334
rect 350 324 351 328
rect 353 330 355 334
rect 359 330 361 334
rect 353 324 361 330
rect 363 328 368 334
rect 586 348 592 363
rect 591 343 592 348
rect 594 347 599 363
rect 594 343 595 347
rect 615 351 621 366
rect 620 346 621 351
rect 623 350 628 366
rect 623 346 624 350
rect 673 348 679 363
rect 678 343 679 348
rect 681 347 686 363
rect 681 343 682 347
rect 702 351 708 366
rect 707 346 708 351
rect 710 350 715 366
rect 710 346 711 350
rect 363 324 364 328
rect 501 315 506 321
rect 290 303 295 309
rect 294 299 295 303
rect 297 305 299 309
rect 303 305 305 309
rect 297 299 305 305
rect 307 303 312 309
rect 307 299 308 303
rect 294 284 295 288
rect 290 268 295 284
rect 297 268 305 288
rect 307 272 312 288
rect 307 268 308 272
rect 195 250 196 254
rect 159 232 164 238
rect 163 228 164 232
rect 166 234 167 238
rect 166 228 171 234
rect 191 214 196 250
rect 198 214 202 254
rect 204 218 209 254
rect 217 250 220 254
rect 213 234 220 250
rect 222 234 229 254
rect 231 238 239 254
rect 243 246 248 252
rect 247 242 248 246
rect 250 248 253 252
rect 467 298 472 314
rect 471 294 472 298
rect 474 294 482 314
rect 484 310 485 314
rect 505 311 506 315
rect 508 317 509 321
rect 508 311 513 317
rect 484 294 489 310
rect 787 331 788 335
rect 751 313 756 319
rect 591 289 596 295
rect 595 285 596 289
rect 598 291 599 295
rect 598 285 603 291
rect 631 285 636 301
rect 635 281 636 285
rect 638 297 639 301
rect 638 281 643 297
rect 755 309 756 313
rect 758 315 759 319
rect 758 309 763 315
rect 678 289 683 295
rect 682 285 683 289
rect 685 291 686 295
rect 685 285 690 291
rect 718 285 723 301
rect 722 281 723 285
rect 725 297 726 301
rect 725 281 730 297
rect 783 295 788 331
rect 790 295 794 335
rect 796 299 801 335
rect 809 331 812 335
rect 805 315 812 331
rect 814 315 821 335
rect 823 319 831 335
rect 835 327 840 333
rect 839 323 840 327
rect 842 329 845 333
rect 842 323 849 329
rect 823 315 827 319
rect 796 295 797 299
rect 250 242 257 248
rect 231 234 235 238
rect 353 235 358 241
rect 357 231 358 235
rect 360 237 362 241
rect 366 237 368 241
rect 360 231 368 237
rect 370 235 375 241
rect 388 239 393 245
rect 392 235 393 239
rect 395 241 396 245
rect 395 235 400 241
rect 370 231 371 235
rect 204 214 205 218
rect 77 139 78 143
rect 41 121 46 127
rect 45 117 46 121
rect 48 123 49 127
rect 48 117 53 123
rect 73 103 78 139
rect 80 103 84 143
rect 86 107 91 143
rect 99 139 102 143
rect 95 123 102 139
rect 104 123 111 143
rect 113 127 121 143
rect 125 135 130 141
rect 129 131 130 135
rect 132 137 135 141
rect 132 131 139 137
rect 428 199 433 215
rect 432 195 433 199
rect 435 195 443 215
rect 445 211 446 215
rect 445 195 450 211
rect 685 216 690 222
rect 473 204 478 210
rect 477 200 478 204
rect 480 206 482 210
rect 486 206 488 210
rect 480 200 488 206
rect 490 204 495 210
rect 508 208 513 214
rect 512 204 513 208
rect 515 210 516 214
rect 689 212 690 216
rect 692 218 693 222
rect 692 212 697 218
rect 787 212 788 216
rect 515 204 520 210
rect 490 200 491 204
rect 670 185 676 200
rect 675 180 676 185
rect 678 184 683 200
rect 678 180 679 184
rect 699 188 705 203
rect 704 183 705 188
rect 707 187 712 203
rect 751 194 756 200
rect 755 190 756 194
rect 758 196 759 200
rect 758 190 763 196
rect 707 183 708 187
rect 603 174 608 180
rect 607 170 608 174
rect 610 176 611 180
rect 783 176 788 212
rect 790 176 794 216
rect 796 180 801 216
rect 809 212 812 216
rect 805 196 812 212
rect 814 196 821 216
rect 823 200 831 216
rect 835 208 840 214
rect 839 204 840 208
rect 842 210 845 214
rect 842 204 849 210
rect 823 196 827 200
rect 796 176 797 180
rect 610 170 615 176
rect 353 137 358 143
rect 357 133 358 137
rect 360 139 362 143
rect 366 139 368 143
rect 360 133 368 139
rect 370 137 375 143
rect 370 133 371 137
rect 588 143 594 158
rect 593 138 594 143
rect 596 142 601 158
rect 596 138 597 142
rect 617 146 623 161
rect 622 141 623 146
rect 625 145 630 161
rect 625 141 626 145
rect 464 131 469 137
rect 113 123 117 127
rect 430 114 435 130
rect 86 103 87 107
rect 292 103 297 109
rect 296 99 297 103
rect 299 105 301 109
rect 305 105 307 109
rect 299 99 307 105
rect 309 103 314 109
rect 309 99 310 103
rect 296 84 297 88
rect 292 68 297 84
rect 299 68 307 88
rect 309 72 314 88
rect 309 68 310 72
rect 434 110 435 114
rect 437 110 445 130
rect 447 126 448 130
rect 468 127 469 131
rect 471 133 472 137
rect 471 127 476 133
rect 447 110 452 126
rect 192 52 193 56
rect 156 34 161 40
rect 160 30 161 34
rect 163 36 164 40
rect 163 30 168 36
rect 188 16 193 52
rect 195 16 199 56
rect 201 20 206 56
rect 214 52 217 56
rect 210 36 217 52
rect 219 36 226 56
rect 228 40 236 56
rect 240 48 245 54
rect 244 44 245 48
rect 247 50 250 54
rect 247 44 254 50
rect 675 126 680 132
rect 679 122 680 126
rect 682 128 683 132
rect 682 122 687 128
rect 715 122 720 138
rect 719 118 720 122
rect 722 134 723 138
rect 722 118 727 134
rect 593 84 598 90
rect 597 80 598 84
rect 600 86 601 90
rect 600 80 605 86
rect 633 80 638 96
rect 637 76 638 80
rect 640 92 641 96
rect 640 76 645 92
rect 790 89 791 93
rect 228 36 232 40
rect 347 47 352 53
rect 351 43 352 47
rect 354 49 356 53
rect 360 49 362 53
rect 354 43 362 49
rect 364 47 369 53
rect 382 51 387 57
rect 386 47 387 51
rect 389 53 390 57
rect 389 47 394 53
rect 754 71 759 77
rect 758 67 759 71
rect 761 73 762 77
rect 761 67 766 73
rect 489 52 494 58
rect 364 43 365 47
rect 406 35 411 51
rect 410 31 411 35
rect 413 31 421 51
rect 423 47 424 51
rect 493 48 494 52
rect 496 54 498 58
rect 502 54 504 58
rect 496 48 504 54
rect 506 52 511 58
rect 524 56 529 62
rect 528 52 529 56
rect 531 58 532 62
rect 531 52 536 58
rect 786 53 791 89
rect 793 53 797 93
rect 799 57 804 93
rect 812 89 815 93
rect 808 73 815 89
rect 817 73 824 93
rect 826 77 834 93
rect 838 85 843 91
rect 842 81 843 85
rect 845 87 848 91
rect 845 81 852 87
rect 826 73 830 77
rect 799 53 800 57
rect 506 48 507 52
rect 423 31 428 47
rect 201 16 202 20
<< pdiffusion >>
rect 182 870 183 874
rect 178 834 183 870
rect 185 834 189 874
rect 191 838 196 874
rect 204 870 205 874
rect 200 854 205 870
rect 207 858 212 874
rect 207 854 208 858
rect 220 870 221 874
rect 216 854 221 870
rect 223 858 228 874
rect 223 854 224 858
rect 266 866 267 870
rect 262 850 267 866
rect 269 854 276 870
rect 269 850 272 854
rect 499 859 500 863
rect 495 843 500 859
rect 502 847 507 863
rect 502 843 503 847
rect 585 857 586 861
rect 191 834 192 838
rect 581 821 586 857
rect 588 821 592 861
rect 594 825 599 861
rect 607 857 608 861
rect 603 841 608 857
rect 610 845 615 861
rect 610 841 611 845
rect 623 857 624 861
rect 619 841 624 857
rect 626 845 631 861
rect 626 841 627 845
rect 669 853 670 857
rect 665 837 670 853
rect 672 841 679 857
rect 672 837 675 841
rect 594 821 595 825
rect 529 775 530 779
rect 337 768 338 772
rect 182 759 183 763
rect 178 723 183 759
rect 185 723 189 763
rect 191 727 196 763
rect 204 759 205 763
rect 200 743 205 759
rect 207 747 212 763
rect 207 743 208 747
rect 220 759 221 763
rect 216 743 221 759
rect 223 747 228 763
rect 223 743 224 747
rect 266 755 267 759
rect 262 739 267 755
rect 269 743 276 759
rect 333 752 338 768
rect 340 756 348 772
rect 340 752 342 756
rect 346 752 348 756
rect 350 768 351 772
rect 350 752 355 768
rect 489 769 490 773
rect 485 753 490 769
rect 492 757 497 773
rect 525 759 530 775
rect 532 763 537 779
rect 532 759 533 763
rect 492 753 493 757
rect 269 739 272 743
rect 681 757 682 761
rect 602 751 603 755
rect 378 736 379 740
rect 191 723 192 727
rect 69 699 70 703
rect 65 663 70 699
rect 72 663 76 703
rect 78 667 83 703
rect 91 699 92 703
rect 87 683 92 699
rect 94 687 99 703
rect 94 683 95 687
rect 107 699 108 703
rect 103 683 108 699
rect 110 687 115 703
rect 110 683 111 687
rect 153 695 154 699
rect 149 679 154 695
rect 156 683 163 699
rect 300 711 301 715
rect 156 679 159 683
rect 296 675 301 711
rect 303 675 311 715
rect 313 679 318 715
rect 374 720 379 736
rect 381 724 386 740
rect 598 735 603 751
rect 605 739 610 755
rect 677 741 682 757
rect 684 745 689 761
rect 684 741 685 745
rect 605 735 606 739
rect 381 720 382 724
rect 743 702 744 706
rect 313 675 314 679
rect 78 663 79 667
rect 369 674 370 678
rect 365 638 370 674
rect 372 638 380 678
rect 382 642 387 678
rect 711 673 712 677
rect 632 667 633 671
rect 592 661 593 665
rect 382 638 383 642
rect 404 654 405 658
rect 400 638 405 654
rect 407 642 412 658
rect 588 645 593 661
rect 595 649 600 665
rect 628 651 633 667
rect 635 655 640 671
rect 635 651 636 655
rect 671 667 672 671
rect 667 651 672 667
rect 674 655 679 671
rect 707 657 712 673
rect 714 661 719 677
rect 739 666 744 702
rect 746 666 750 706
rect 752 670 757 706
rect 765 702 766 706
rect 761 686 766 702
rect 768 690 773 706
rect 768 686 769 690
rect 781 702 782 706
rect 777 686 782 702
rect 784 690 789 706
rect 784 686 785 690
rect 827 698 828 702
rect 823 682 828 698
rect 830 686 837 702
rect 830 682 833 686
rect 752 666 753 670
rect 714 657 715 661
rect 674 651 675 655
rect 595 645 596 649
rect 407 638 408 642
rect 172 620 173 624
rect 168 584 173 620
rect 175 584 179 624
rect 181 588 186 624
rect 194 620 195 624
rect 190 604 195 620
rect 197 608 202 624
rect 197 604 198 608
rect 210 620 211 624
rect 206 604 211 620
rect 213 608 218 624
rect 213 604 214 608
rect 256 616 257 620
rect 252 600 257 616
rect 259 604 266 620
rect 435 629 436 633
rect 259 600 262 604
rect 431 613 436 629
rect 438 617 446 633
rect 438 613 440 617
rect 444 613 446 617
rect 448 629 449 633
rect 448 613 453 629
rect 181 584 182 588
rect 61 558 62 562
rect 57 522 62 558
rect 64 522 68 562
rect 70 526 75 562
rect 83 558 84 562
rect 79 542 84 558
rect 86 546 91 562
rect 86 542 87 546
rect 99 558 100 562
rect 95 542 100 558
rect 102 546 107 562
rect 102 542 103 546
rect 145 554 146 558
rect 141 538 146 554
rect 148 542 155 558
rect 296 579 301 595
rect 300 575 301 579
rect 303 591 305 595
rect 309 591 311 595
rect 303 575 311 591
rect 313 579 318 595
rect 313 575 314 579
rect 369 576 370 580
rect 148 538 151 542
rect 70 522 71 526
rect 295 537 296 541
rect 291 501 296 537
rect 298 501 306 541
rect 308 505 313 541
rect 365 540 370 576
rect 372 540 380 580
rect 382 544 387 580
rect 600 579 601 583
rect 596 563 601 579
rect 603 567 608 583
rect 603 563 604 567
rect 691 579 692 583
rect 687 563 692 579
rect 694 567 699 583
rect 694 563 695 567
rect 382 540 383 544
rect 427 544 428 548
rect 423 528 428 544
rect 430 532 438 548
rect 430 528 432 532
rect 436 528 438 532
rect 440 544 441 548
rect 440 528 445 544
rect 461 544 462 548
rect 457 528 462 544
rect 464 532 469 548
rect 464 528 465 532
rect 308 501 309 505
rect 359 486 360 490
rect 170 459 171 463
rect 166 423 171 459
rect 173 423 177 463
rect 179 427 184 463
rect 192 459 193 463
rect 188 443 193 459
rect 195 447 200 463
rect 195 443 196 447
rect 208 459 209 463
rect 204 443 209 459
rect 211 447 216 463
rect 211 443 212 447
rect 254 455 255 459
rect 250 439 255 455
rect 257 443 264 459
rect 257 439 260 443
rect 355 450 360 486
rect 362 450 370 490
rect 372 454 377 490
rect 755 524 756 528
rect 630 495 631 499
rect 590 489 591 493
rect 482 481 483 485
rect 372 450 373 454
rect 394 466 395 470
rect 390 450 395 466
rect 397 454 402 470
rect 397 450 398 454
rect 179 423 180 427
rect 46 405 47 409
rect 42 369 47 405
rect 49 369 53 409
rect 55 373 60 409
rect 68 405 69 409
rect 64 389 69 405
rect 71 393 76 409
rect 71 389 72 393
rect 84 405 85 409
rect 80 389 85 405
rect 87 393 92 409
rect 87 389 88 393
rect 130 401 131 405
rect 126 385 131 401
rect 133 389 140 405
rect 133 385 136 389
rect 432 442 433 446
rect 428 426 433 442
rect 435 430 443 446
rect 435 426 437 430
rect 441 426 443 430
rect 445 442 446 446
rect 478 445 483 481
rect 485 445 493 485
rect 495 449 500 485
rect 586 473 591 489
rect 593 477 598 493
rect 626 479 631 495
rect 633 483 638 499
rect 721 495 722 499
rect 633 479 634 483
rect 681 489 682 493
rect 593 473 594 477
rect 495 445 496 449
rect 517 461 518 465
rect 513 445 518 461
rect 520 449 525 465
rect 677 473 682 489
rect 684 477 689 493
rect 717 479 722 495
rect 724 483 729 499
rect 751 488 756 524
rect 758 488 762 528
rect 764 492 769 528
rect 777 524 778 528
rect 773 508 778 524
rect 780 512 785 528
rect 780 508 781 512
rect 793 524 794 528
rect 789 508 794 524
rect 796 512 801 528
rect 796 508 797 512
rect 839 520 840 524
rect 835 504 840 520
rect 842 508 849 524
rect 842 504 845 508
rect 764 488 765 492
rect 724 479 725 483
rect 684 473 685 477
rect 520 445 521 449
rect 445 426 450 442
rect 291 405 296 421
rect 295 401 296 405
rect 298 417 300 421
rect 304 417 306 421
rect 298 401 306 417
rect 308 405 313 421
rect 605 413 606 417
rect 308 401 309 405
rect 350 388 351 392
rect 55 369 56 373
rect 294 364 295 368
rect 290 328 295 364
rect 297 328 305 368
rect 307 332 312 368
rect 346 352 351 388
rect 353 352 361 392
rect 363 356 368 392
rect 601 397 606 413
rect 608 401 613 417
rect 608 397 609 401
rect 692 413 693 417
rect 688 397 693 413
rect 695 401 700 417
rect 695 397 696 401
rect 363 352 364 356
rect 471 349 472 353
rect 307 328 308 332
rect 467 333 472 349
rect 474 337 482 353
rect 474 333 476 337
rect 480 333 482 337
rect 484 349 485 353
rect 484 333 489 349
rect 505 349 506 353
rect 501 333 506 349
rect 508 337 513 353
rect 755 367 756 371
rect 508 333 509 337
rect 635 329 636 333
rect 595 323 596 327
rect 357 295 358 299
rect 163 286 164 290
rect 159 250 164 286
rect 166 250 170 290
rect 172 254 177 290
rect 185 286 186 290
rect 181 270 186 286
rect 188 274 193 290
rect 188 270 189 274
rect 201 286 202 290
rect 197 270 202 286
rect 204 274 209 290
rect 204 270 205 274
rect 247 282 248 286
rect 243 266 248 282
rect 250 270 257 286
rect 250 266 253 270
rect 172 250 173 254
rect 353 259 358 295
rect 360 259 368 299
rect 370 263 375 299
rect 591 307 596 323
rect 598 311 603 327
rect 631 313 636 329
rect 638 317 643 333
rect 722 329 723 333
rect 638 313 639 317
rect 682 323 683 327
rect 598 307 599 311
rect 678 307 683 323
rect 685 311 690 327
rect 718 313 723 329
rect 725 317 730 333
rect 751 331 756 367
rect 758 331 762 371
rect 764 335 769 371
rect 777 367 778 371
rect 773 351 778 367
rect 780 355 785 371
rect 780 351 781 355
rect 793 367 794 371
rect 789 351 794 367
rect 796 355 801 371
rect 796 351 797 355
rect 839 363 840 367
rect 835 347 840 363
rect 842 351 849 367
rect 842 347 845 351
rect 764 331 765 335
rect 725 313 726 317
rect 685 307 686 311
rect 370 259 371 263
rect 392 275 393 279
rect 388 259 393 275
rect 395 263 400 279
rect 395 259 396 263
rect 477 264 478 268
rect 290 232 295 248
rect 294 228 295 232
rect 297 244 299 248
rect 303 244 305 248
rect 297 228 305 244
rect 307 232 312 248
rect 432 250 433 254
rect 307 228 308 232
rect 428 234 433 250
rect 435 238 443 254
rect 435 234 437 238
rect 441 234 443 238
rect 445 250 446 254
rect 445 234 450 250
rect 473 228 478 264
rect 480 228 488 268
rect 490 232 495 268
rect 689 250 690 254
rect 490 228 491 232
rect 512 244 513 248
rect 508 228 513 244
rect 515 232 520 248
rect 685 234 690 250
rect 692 238 697 254
rect 692 234 693 238
rect 755 248 756 252
rect 515 228 516 232
rect 357 197 358 201
rect 45 175 46 179
rect 41 139 46 175
rect 48 139 52 179
rect 54 143 59 179
rect 67 175 68 179
rect 63 159 68 175
rect 70 163 75 179
rect 70 159 71 163
rect 83 175 84 179
rect 79 159 84 175
rect 86 163 91 179
rect 86 159 87 163
rect 129 171 130 175
rect 125 155 130 171
rect 132 159 139 175
rect 132 155 135 159
rect 296 164 297 168
rect 54 139 55 143
rect 292 128 297 164
rect 299 128 307 168
rect 309 132 314 168
rect 353 161 358 197
rect 360 161 368 201
rect 370 165 375 201
rect 751 212 756 248
rect 758 212 762 252
rect 764 216 769 252
rect 777 248 778 252
rect 773 232 778 248
rect 780 236 785 252
rect 780 232 781 236
rect 793 248 794 252
rect 789 232 794 248
rect 796 236 801 252
rect 796 232 797 236
rect 839 244 840 248
rect 835 228 840 244
rect 842 232 849 248
rect 842 228 845 232
rect 764 212 765 216
rect 607 208 608 212
rect 603 192 608 208
rect 610 196 615 212
rect 610 192 611 196
rect 370 161 371 165
rect 434 165 435 169
rect 430 149 435 165
rect 437 153 445 169
rect 437 149 439 153
rect 443 149 445 153
rect 447 165 448 169
rect 447 149 452 165
rect 468 165 469 169
rect 464 149 469 165
rect 471 153 476 169
rect 719 166 720 170
rect 471 149 472 153
rect 309 128 310 132
rect 679 160 680 164
rect 675 144 680 160
rect 682 148 687 164
rect 715 150 720 166
rect 722 154 727 170
rect 722 150 723 154
rect 682 144 683 148
rect 351 107 352 111
rect 160 88 161 92
rect 156 52 161 88
rect 163 52 167 92
rect 169 56 174 92
rect 182 88 183 92
rect 178 72 183 88
rect 185 76 190 92
rect 185 72 186 76
rect 198 88 199 92
rect 194 72 199 88
rect 201 76 206 92
rect 201 72 202 76
rect 244 84 245 88
rect 240 68 245 84
rect 247 72 254 88
rect 247 68 250 72
rect 347 71 352 107
rect 354 71 362 111
rect 364 75 369 111
rect 637 124 638 128
rect 597 118 598 122
rect 493 112 494 116
rect 364 71 365 75
rect 386 87 387 91
rect 382 71 387 87
rect 389 75 394 91
rect 389 71 390 75
rect 410 86 411 90
rect 169 52 170 56
rect 406 70 411 86
rect 413 74 421 90
rect 413 70 415 74
rect 419 70 421 74
rect 423 86 424 90
rect 423 70 428 86
rect 489 76 494 112
rect 496 76 504 116
rect 506 80 511 116
rect 593 102 598 118
rect 600 106 605 122
rect 633 108 638 124
rect 640 112 645 128
rect 758 125 759 129
rect 640 108 641 112
rect 600 102 601 106
rect 506 76 507 80
rect 528 92 529 96
rect 524 76 529 92
rect 531 80 536 96
rect 531 76 532 80
rect 754 89 759 125
rect 761 89 765 129
rect 767 93 772 129
rect 780 125 781 129
rect 776 109 781 125
rect 783 113 788 129
rect 783 109 784 113
rect 796 125 797 129
rect 792 109 797 125
rect 799 113 804 129
rect 799 109 800 113
rect 842 121 843 125
rect 838 105 843 121
rect 845 109 852 125
rect 845 105 848 109
rect 767 89 768 93
rect 292 32 297 48
rect 296 28 297 32
rect 299 44 301 48
rect 305 44 307 48
rect 299 28 307 44
rect 309 32 314 48
rect 309 28 310 32
<< ndcontact >>
rect 210 834 214 838
rect 178 812 182 816
rect 186 818 190 822
rect 232 834 236 838
rect 262 826 266 830
rect 272 832 276 836
rect 254 818 258 822
rect 495 821 499 825
rect 503 827 507 831
rect 613 821 617 825
rect 224 798 228 802
rect 489 789 493 793
rect 581 799 585 803
rect 589 805 593 809
rect 518 792 522 796
rect 635 821 639 825
rect 665 813 669 817
rect 675 819 679 823
rect 657 805 661 809
rect 627 785 631 789
rect 210 723 214 727
rect 178 701 182 705
rect 186 707 190 711
rect 232 723 236 727
rect 262 715 266 719
rect 272 721 276 725
rect 254 707 258 711
rect 224 687 228 691
rect 333 713 337 717
rect 351 729 355 733
rect 485 731 489 735
rect 493 737 497 741
rect 525 727 529 731
rect 533 743 537 747
rect 598 713 602 717
rect 606 719 610 723
rect 677 719 681 723
rect 685 725 689 729
rect 374 698 378 702
rect 382 704 386 708
rect 592 681 596 685
rect 621 684 625 688
rect 671 687 675 691
rect 700 690 704 694
rect 97 663 101 667
rect 65 641 69 645
rect 73 647 77 651
rect 119 663 123 667
rect 149 655 153 659
rect 159 661 163 665
rect 141 647 145 651
rect 296 646 300 650
rect 305 652 309 656
rect 314 646 318 650
rect 771 666 775 670
rect 111 627 115 631
rect 296 631 300 635
rect 314 615 318 619
rect 365 610 369 614
rect 374 616 378 620
rect 400 614 404 618
rect 408 620 412 624
rect 383 610 387 614
rect 588 623 592 627
rect 596 629 600 633
rect 628 619 632 623
rect 636 635 640 639
rect 667 629 671 633
rect 675 635 679 639
rect 707 625 711 629
rect 715 641 719 645
rect 739 644 743 648
rect 747 650 751 654
rect 793 666 797 670
rect 823 658 827 662
rect 833 664 837 668
rect 815 650 819 654
rect 785 630 789 634
rect 200 584 204 588
rect 168 562 172 566
rect 176 568 180 572
rect 222 584 226 588
rect 252 576 256 580
rect 262 582 266 586
rect 244 568 248 572
rect 214 548 218 552
rect 89 522 93 526
rect 57 500 61 504
rect 65 506 69 510
rect 111 522 115 526
rect 141 514 145 518
rect 151 520 155 524
rect 133 506 137 510
rect 431 574 435 578
rect 449 590 453 594
rect 596 541 600 545
rect 604 547 608 551
rect 687 541 691 545
rect 695 547 699 551
rect 365 512 369 516
rect 374 518 378 522
rect 383 512 387 516
rect 103 486 107 490
rect 291 472 295 476
rect 300 478 304 482
rect 309 472 313 476
rect 291 457 295 461
rect 423 489 427 493
rect 441 505 445 509
rect 457 506 461 510
rect 465 512 469 516
rect 590 509 594 513
rect 619 512 623 516
rect 681 509 685 513
rect 710 512 714 516
rect 309 441 313 445
rect 198 423 202 427
rect 166 401 170 405
rect 174 407 178 411
rect 220 423 224 427
rect 250 415 254 419
rect 260 421 264 425
rect 355 422 359 426
rect 364 428 368 432
rect 390 426 394 430
rect 398 432 402 436
rect 783 488 787 492
rect 586 451 590 455
rect 594 457 598 461
rect 626 447 630 451
rect 634 463 638 467
rect 677 451 681 455
rect 685 457 689 461
rect 717 447 721 451
rect 725 463 729 467
rect 751 466 755 470
rect 759 472 763 476
rect 805 488 809 492
rect 835 480 839 484
rect 845 486 849 490
rect 827 472 831 476
rect 797 452 801 456
rect 373 422 377 426
rect 242 407 246 411
rect 478 417 482 421
rect 487 423 491 427
rect 513 421 517 425
rect 521 427 525 431
rect 496 417 500 421
rect 212 387 216 391
rect 74 369 78 373
rect 42 347 46 351
rect 50 353 54 357
rect 96 369 100 373
rect 126 361 130 365
rect 136 367 140 371
rect 118 353 122 357
rect 88 333 92 337
rect 428 387 432 391
rect 446 403 450 407
rect 601 375 605 379
rect 609 381 613 385
rect 688 375 692 379
rect 696 381 700 385
rect 346 324 350 328
rect 355 330 359 334
rect 595 343 599 347
rect 624 346 628 350
rect 682 343 686 347
rect 711 346 715 350
rect 364 324 368 328
rect 290 299 294 303
rect 299 305 303 309
rect 308 299 312 303
rect 290 284 294 288
rect 308 268 312 272
rect 191 250 195 254
rect 159 228 163 232
rect 167 234 171 238
rect 213 250 217 254
rect 243 242 247 246
rect 253 248 257 252
rect 467 294 471 298
rect 485 310 489 314
rect 501 311 505 315
rect 509 317 513 321
rect 783 331 787 335
rect 591 285 595 289
rect 599 291 603 295
rect 631 281 635 285
rect 639 297 643 301
rect 751 309 755 313
rect 759 315 763 319
rect 678 285 682 289
rect 686 291 690 295
rect 718 281 722 285
rect 726 297 730 301
rect 805 331 809 335
rect 835 323 839 327
rect 845 329 849 333
rect 827 315 831 319
rect 797 295 801 299
rect 235 234 239 238
rect 353 231 357 235
rect 362 237 366 241
rect 388 235 392 239
rect 396 241 400 245
rect 371 231 375 235
rect 205 214 209 218
rect 73 139 77 143
rect 41 117 45 121
rect 49 123 53 127
rect 95 139 99 143
rect 125 131 129 135
rect 135 137 139 141
rect 428 195 432 199
rect 446 211 450 215
rect 473 200 477 204
rect 482 206 486 210
rect 508 204 512 208
rect 516 210 520 214
rect 685 212 689 216
rect 693 218 697 222
rect 783 212 787 216
rect 491 200 495 204
rect 679 180 683 184
rect 751 190 755 194
rect 759 196 763 200
rect 708 183 712 187
rect 603 170 607 174
rect 611 176 615 180
rect 805 212 809 216
rect 835 204 839 208
rect 845 210 849 214
rect 827 196 831 200
rect 797 176 801 180
rect 353 133 357 137
rect 362 139 366 143
rect 371 133 375 137
rect 597 138 601 142
rect 626 141 630 145
rect 117 123 121 127
rect 87 103 91 107
rect 292 99 296 103
rect 301 105 305 109
rect 310 99 314 103
rect 292 84 296 88
rect 310 68 314 72
rect 430 110 434 114
rect 448 126 452 130
rect 464 127 468 131
rect 472 133 476 137
rect 188 52 192 56
rect 156 30 160 34
rect 164 36 168 40
rect 210 52 214 56
rect 240 44 244 48
rect 250 50 254 54
rect 675 122 679 126
rect 683 128 687 132
rect 715 118 719 122
rect 723 134 727 138
rect 593 80 597 84
rect 601 86 605 90
rect 633 76 637 80
rect 641 92 645 96
rect 786 89 790 93
rect 232 36 236 40
rect 347 43 351 47
rect 356 49 360 53
rect 382 47 386 51
rect 390 53 394 57
rect 754 67 758 71
rect 762 73 766 77
rect 365 43 369 47
rect 406 31 410 35
rect 424 47 428 51
rect 489 48 493 52
rect 498 54 502 58
rect 524 52 528 56
rect 532 58 536 62
rect 808 89 812 93
rect 838 81 842 85
rect 848 87 852 91
rect 830 73 834 77
rect 800 53 804 57
rect 507 48 511 52
rect 202 16 206 20
<< pdcontact >>
rect 178 870 182 874
rect 200 870 204 874
rect 208 854 212 858
rect 216 870 220 874
rect 224 854 228 858
rect 262 866 266 870
rect 272 850 276 854
rect 495 859 499 863
rect 503 843 507 847
rect 581 857 585 861
rect 192 834 196 838
rect 603 857 607 861
rect 611 841 615 845
rect 619 857 623 861
rect 627 841 631 845
rect 665 853 669 857
rect 675 837 679 841
rect 595 821 599 825
rect 525 775 529 779
rect 333 768 337 772
rect 178 759 182 763
rect 200 759 204 763
rect 208 743 212 747
rect 216 759 220 763
rect 224 743 228 747
rect 262 755 266 759
rect 342 752 346 756
rect 351 768 355 772
rect 485 769 489 773
rect 533 759 537 763
rect 493 753 497 757
rect 272 739 276 743
rect 677 757 681 761
rect 598 751 602 755
rect 374 736 378 740
rect 192 723 196 727
rect 65 699 69 703
rect 87 699 91 703
rect 95 683 99 687
rect 103 699 107 703
rect 111 683 115 687
rect 149 695 153 699
rect 296 711 300 715
rect 159 679 163 683
rect 685 741 689 745
rect 606 735 610 739
rect 382 720 386 724
rect 739 702 743 706
rect 314 675 318 679
rect 79 663 83 667
rect 365 674 369 678
rect 707 673 711 677
rect 628 667 632 671
rect 588 661 592 665
rect 383 638 387 642
rect 400 654 404 658
rect 636 651 640 655
rect 667 667 671 671
rect 761 702 765 706
rect 769 686 773 690
rect 777 702 781 706
rect 785 686 789 690
rect 823 698 827 702
rect 833 682 837 686
rect 753 666 757 670
rect 715 657 719 661
rect 675 651 679 655
rect 596 645 600 649
rect 408 638 412 642
rect 168 620 172 624
rect 190 620 194 624
rect 198 604 202 608
rect 206 620 210 624
rect 214 604 218 608
rect 252 616 256 620
rect 431 629 435 633
rect 262 600 266 604
rect 440 613 444 617
rect 449 629 453 633
rect 182 584 186 588
rect 57 558 61 562
rect 79 558 83 562
rect 87 542 91 546
rect 95 558 99 562
rect 103 542 107 546
rect 141 554 145 558
rect 296 575 300 579
rect 305 591 309 595
rect 314 575 318 579
rect 365 576 369 580
rect 151 538 155 542
rect 71 522 75 526
rect 291 537 295 541
rect 596 579 600 583
rect 604 563 608 567
rect 687 579 691 583
rect 695 563 699 567
rect 383 540 387 544
rect 423 544 427 548
rect 432 528 436 532
rect 441 544 445 548
rect 457 544 461 548
rect 465 528 469 532
rect 309 501 313 505
rect 355 486 359 490
rect 166 459 170 463
rect 188 459 192 463
rect 196 443 200 447
rect 204 459 208 463
rect 212 443 216 447
rect 250 455 254 459
rect 260 439 264 443
rect 751 524 755 528
rect 626 495 630 499
rect 586 489 590 493
rect 478 481 482 485
rect 373 450 377 454
rect 390 466 394 470
rect 398 450 402 454
rect 180 423 184 427
rect 42 405 46 409
rect 64 405 68 409
rect 72 389 76 393
rect 80 405 84 409
rect 88 389 92 393
rect 126 401 130 405
rect 136 385 140 389
rect 428 442 432 446
rect 437 426 441 430
rect 446 442 450 446
rect 717 495 721 499
rect 634 479 638 483
rect 677 489 681 493
rect 594 473 598 477
rect 496 445 500 449
rect 513 461 517 465
rect 773 524 777 528
rect 781 508 785 512
rect 789 524 793 528
rect 797 508 801 512
rect 835 520 839 524
rect 845 504 849 508
rect 765 488 769 492
rect 725 479 729 483
rect 685 473 689 477
rect 521 445 525 449
rect 291 401 295 405
rect 300 417 304 421
rect 601 413 605 417
rect 309 401 313 405
rect 346 388 350 392
rect 56 369 60 373
rect 290 364 294 368
rect 609 397 613 401
rect 688 413 692 417
rect 696 397 700 401
rect 364 352 368 356
rect 467 349 471 353
rect 308 328 312 332
rect 476 333 480 337
rect 485 349 489 353
rect 501 349 505 353
rect 751 367 755 371
rect 509 333 513 337
rect 631 329 635 333
rect 591 323 595 327
rect 353 295 357 299
rect 159 286 163 290
rect 181 286 185 290
rect 189 270 193 274
rect 197 286 201 290
rect 205 270 209 274
rect 243 282 247 286
rect 253 266 257 270
rect 173 250 177 254
rect 718 329 722 333
rect 639 313 643 317
rect 678 323 682 327
rect 599 307 603 311
rect 773 367 777 371
rect 781 351 785 355
rect 789 367 793 371
rect 797 351 801 355
rect 835 363 839 367
rect 845 347 849 351
rect 765 331 769 335
rect 726 313 730 317
rect 686 307 690 311
rect 371 259 375 263
rect 388 275 392 279
rect 396 259 400 263
rect 473 264 477 268
rect 290 228 294 232
rect 299 244 303 248
rect 428 250 432 254
rect 308 228 312 232
rect 437 234 441 238
rect 446 250 450 254
rect 685 250 689 254
rect 491 228 495 232
rect 508 244 512 248
rect 693 234 697 238
rect 751 248 755 252
rect 516 228 520 232
rect 353 197 357 201
rect 41 175 45 179
rect 63 175 67 179
rect 71 159 75 163
rect 79 175 83 179
rect 87 159 91 163
rect 125 171 129 175
rect 135 155 139 159
rect 292 164 296 168
rect 55 139 59 143
rect 773 248 777 252
rect 781 232 785 236
rect 789 248 793 252
rect 797 232 801 236
rect 835 244 839 248
rect 845 228 849 232
rect 765 212 769 216
rect 603 208 607 212
rect 611 192 615 196
rect 371 161 375 165
rect 430 165 434 169
rect 439 149 443 153
rect 448 165 452 169
rect 464 165 468 169
rect 715 166 719 170
rect 472 149 476 153
rect 310 128 314 132
rect 675 160 679 164
rect 723 150 727 154
rect 683 144 687 148
rect 347 107 351 111
rect 156 88 160 92
rect 178 88 182 92
rect 186 72 190 76
rect 194 88 198 92
rect 202 72 206 76
rect 240 84 244 88
rect 250 68 254 72
rect 633 124 637 128
rect 593 118 597 122
rect 489 112 493 116
rect 365 71 369 75
rect 382 87 386 91
rect 390 71 394 75
rect 406 86 410 90
rect 170 52 174 56
rect 415 70 419 74
rect 424 86 428 90
rect 754 125 758 129
rect 641 108 645 112
rect 601 102 605 106
rect 507 76 511 80
rect 524 92 528 96
rect 532 76 536 80
rect 776 125 780 129
rect 784 109 788 113
rect 792 125 796 129
rect 800 109 804 113
rect 838 121 842 125
rect 848 105 852 109
rect 768 89 772 93
rect 292 28 296 32
rect 301 44 305 48
rect 310 28 314 32
<< polysilicon >>
rect 183 874 185 877
rect 189 874 191 881
rect 205 874 207 886
rect 221 874 223 877
rect 267 870 269 878
rect 205 851 207 854
rect 221 849 223 854
rect 500 863 502 866
rect 215 838 217 841
rect 267 843 269 850
rect 586 861 588 864
rect 592 861 594 868
rect 608 861 610 873
rect 624 861 626 864
rect 221 838 223 839
rect 239 838 241 839
rect 248 838 250 841
rect 183 822 185 834
rect 189 831 191 834
rect 183 809 185 812
rect 267 836 269 839
rect 500 831 502 843
rect 267 823 269 826
rect 670 857 672 865
rect 608 838 610 841
rect 624 836 626 841
rect 618 825 620 828
rect 670 830 672 837
rect 624 825 626 826
rect 642 825 644 826
rect 651 825 653 828
rect 500 818 502 821
rect 239 815 241 818
rect 248 815 250 818
rect 515 812 517 813
rect 486 809 488 810
rect 215 797 217 798
rect 221 795 223 798
rect 586 809 588 821
rect 592 818 594 821
rect 586 796 588 799
rect 515 789 517 792
rect 486 786 488 789
rect 670 823 672 826
rect 670 810 672 813
rect 642 802 644 805
rect 651 802 653 805
rect 618 784 620 785
rect 530 779 532 782
rect 624 782 626 785
rect 183 763 185 766
rect 189 763 191 770
rect 205 763 207 775
rect 338 772 340 776
rect 348 772 350 776
rect 490 773 492 776
rect 221 763 223 766
rect 267 759 269 767
rect 205 740 207 743
rect 221 738 223 743
rect 682 761 684 764
rect 215 727 217 730
rect 267 732 269 739
rect 338 733 340 752
rect 348 733 350 752
rect 379 740 381 743
rect 490 741 492 753
rect 530 747 532 759
rect 603 755 605 758
rect 221 727 223 728
rect 239 727 241 728
rect 248 727 250 730
rect 70 703 72 706
rect 76 703 78 710
rect 92 703 94 715
rect 183 711 185 723
rect 189 720 191 723
rect 108 703 110 706
rect 154 699 156 707
rect 92 680 94 683
rect 108 678 110 683
rect 183 698 185 701
rect 267 725 269 728
rect 301 715 303 718
rect 311 715 313 718
rect 267 712 269 715
rect 239 704 241 707
rect 248 704 250 707
rect 215 686 217 687
rect 221 684 223 687
rect 102 667 104 670
rect 154 672 156 679
rect 490 728 492 731
rect 530 724 532 727
rect 603 723 605 735
rect 682 729 684 741
rect 338 710 340 713
rect 348 710 350 713
rect 379 708 381 720
rect 682 716 684 719
rect 603 710 605 713
rect 697 710 699 711
rect 668 707 670 708
rect 618 704 620 705
rect 589 701 591 702
rect 379 695 381 698
rect 744 706 746 709
rect 750 706 752 713
rect 766 706 768 718
rect 782 706 784 709
rect 697 687 699 690
rect 668 684 670 687
rect 618 681 620 684
rect 370 678 372 681
rect 380 678 382 681
rect 589 678 591 681
rect 108 667 110 668
rect 126 667 128 668
rect 135 667 137 670
rect 70 651 72 663
rect 76 660 78 663
rect 70 638 72 641
rect 154 665 156 668
rect 301 656 303 675
rect 311 656 313 675
rect 154 652 156 655
rect 126 644 128 647
rect 135 644 137 647
rect 301 643 303 646
rect 311 643 313 646
rect 712 677 714 680
rect 633 671 635 674
rect 672 671 674 674
rect 593 665 595 668
rect 405 658 407 661
rect 828 702 830 710
rect 766 683 768 686
rect 782 681 784 686
rect 776 670 778 673
rect 828 675 830 682
rect 782 670 784 671
rect 800 670 802 671
rect 809 670 811 673
rect 102 626 104 627
rect 108 624 110 627
rect 173 624 175 627
rect 179 624 181 631
rect 195 624 197 636
rect 301 635 303 638
rect 311 635 313 638
rect 211 624 213 627
rect 257 620 259 628
rect 195 601 197 604
rect 211 599 213 604
rect 370 620 372 638
rect 380 620 382 638
rect 405 624 407 638
rect 436 633 438 637
rect 446 633 448 637
rect 593 633 595 645
rect 633 639 635 651
rect 672 639 674 651
rect 712 645 714 657
rect 744 654 746 666
rect 750 663 752 666
rect 205 588 207 591
rect 257 593 259 600
rect 301 595 303 615
rect 311 595 313 615
rect 405 611 407 614
rect 593 620 595 623
rect 672 626 674 629
rect 744 641 746 644
rect 828 668 830 671
rect 828 655 830 658
rect 800 647 802 650
rect 809 647 811 650
rect 776 629 778 630
rect 782 627 784 630
rect 712 622 714 625
rect 633 616 635 619
rect 370 607 372 610
rect 380 607 382 610
rect 211 588 213 589
rect 229 588 231 589
rect 238 588 240 591
rect 62 562 64 565
rect 68 562 70 569
rect 84 562 86 574
rect 173 572 175 584
rect 179 581 181 584
rect 100 562 102 565
rect 146 558 148 566
rect 173 559 175 562
rect 84 539 86 542
rect 100 537 102 542
rect 257 586 259 589
rect 257 573 259 576
rect 436 594 438 613
rect 446 594 448 613
rect 370 580 372 583
rect 380 580 382 583
rect 301 571 303 575
rect 311 571 313 575
rect 229 565 231 568
rect 238 565 240 568
rect 205 547 207 548
rect 211 545 213 548
rect 296 541 298 544
rect 306 541 308 544
rect 94 526 96 529
rect 146 531 148 538
rect 100 526 102 527
rect 118 526 120 527
rect 127 526 129 529
rect 62 510 64 522
rect 68 519 70 522
rect 62 497 64 500
rect 146 524 148 527
rect 146 511 148 514
rect 118 503 120 506
rect 127 503 129 506
rect 601 583 603 586
rect 692 583 694 586
rect 436 571 438 574
rect 446 571 448 574
rect 428 548 430 552
rect 438 548 440 552
rect 601 551 603 563
rect 692 551 694 563
rect 462 548 464 551
rect 370 522 372 540
rect 380 522 382 540
rect 601 538 603 541
rect 692 538 694 541
rect 616 532 618 533
rect 587 529 589 530
rect 370 509 372 512
rect 380 509 382 512
rect 428 509 430 528
rect 438 509 440 528
rect 462 516 464 528
rect 94 485 96 486
rect 100 483 102 486
rect 296 482 298 501
rect 306 482 308 501
rect 360 490 362 493
rect 370 490 372 493
rect 171 463 173 466
rect 177 463 179 470
rect 193 463 195 475
rect 296 469 298 472
rect 306 469 308 472
rect 209 463 211 466
rect 255 459 257 467
rect 296 461 298 464
rect 306 461 308 464
rect 193 440 195 443
rect 209 438 211 443
rect 707 532 709 533
rect 678 529 680 530
rect 616 509 618 512
rect 756 528 758 531
rect 762 528 764 535
rect 778 528 780 540
rect 794 528 796 531
rect 707 509 709 512
rect 587 506 589 509
rect 678 506 680 509
rect 462 503 464 506
rect 631 499 633 502
rect 722 499 724 502
rect 591 493 593 496
rect 428 486 430 489
rect 438 486 440 489
rect 483 485 485 488
rect 493 485 495 488
rect 395 470 397 473
rect 203 427 205 430
rect 255 432 257 439
rect 209 427 211 428
rect 227 427 229 428
rect 236 427 238 430
rect 47 409 49 412
rect 53 409 55 416
rect 69 409 71 421
rect 85 409 87 412
rect 131 405 133 413
rect 171 411 173 423
rect 177 420 179 423
rect 69 386 71 389
rect 85 384 87 389
rect 171 398 173 401
rect 255 425 257 428
rect 296 421 298 441
rect 306 421 308 441
rect 360 432 362 450
rect 370 432 372 450
rect 395 436 397 450
rect 433 446 435 450
rect 443 446 445 450
rect 682 493 684 496
rect 518 465 520 468
rect 591 461 593 473
rect 631 467 633 479
rect 840 524 842 532
rect 778 505 780 508
rect 794 503 796 508
rect 788 492 790 495
rect 840 497 842 504
rect 794 492 796 493
rect 812 492 814 493
rect 821 492 823 495
rect 591 448 593 451
rect 682 461 684 473
rect 722 467 724 479
rect 756 476 758 488
rect 762 485 764 488
rect 682 448 684 451
rect 756 463 758 466
rect 840 490 842 493
rect 840 477 842 480
rect 812 469 814 472
rect 821 469 823 472
rect 788 451 790 452
rect 794 449 796 452
rect 483 427 485 445
rect 493 427 495 445
rect 518 431 520 445
rect 631 444 633 447
rect 722 444 724 447
rect 395 423 397 426
rect 255 412 257 415
rect 227 404 229 407
rect 236 404 238 407
rect 360 419 362 422
rect 370 419 372 422
rect 433 407 435 426
rect 443 407 445 426
rect 518 418 520 421
rect 606 417 608 420
rect 693 417 695 420
rect 483 414 485 417
rect 493 414 495 417
rect 296 397 298 401
rect 306 397 308 401
rect 351 392 353 395
rect 361 392 363 395
rect 203 386 205 387
rect 79 373 81 376
rect 131 378 133 385
rect 209 384 211 387
rect 85 373 87 374
rect 103 373 105 374
rect 112 373 114 376
rect 47 357 49 369
rect 53 366 55 369
rect 47 344 49 347
rect 131 371 133 374
rect 295 368 297 371
rect 305 368 307 371
rect 131 358 133 361
rect 103 350 105 353
rect 112 350 114 353
rect 79 332 81 333
rect 85 330 87 333
rect 433 384 435 387
rect 443 384 445 387
rect 606 385 608 397
rect 693 385 695 397
rect 606 372 608 375
rect 693 372 695 375
rect 756 371 758 374
rect 762 371 764 378
rect 778 371 780 383
rect 794 371 796 374
rect 621 366 623 367
rect 592 363 594 364
rect 472 353 474 357
rect 482 353 484 357
rect 506 353 508 356
rect 351 334 353 352
rect 361 334 363 352
rect 295 309 297 328
rect 305 309 307 328
rect 708 366 710 367
rect 679 363 681 364
rect 621 343 623 346
rect 708 343 710 346
rect 592 340 594 343
rect 679 340 681 343
rect 636 333 638 336
rect 723 333 725 336
rect 351 321 353 324
rect 361 321 363 324
rect 472 314 474 333
rect 482 314 484 333
rect 506 321 508 333
rect 596 327 598 330
rect 164 290 166 293
rect 170 290 172 297
rect 186 290 188 302
rect 358 299 360 302
rect 368 299 370 302
rect 295 296 297 299
rect 305 296 307 299
rect 202 290 204 293
rect 248 286 250 294
rect 295 288 297 291
rect 305 288 307 291
rect 186 267 188 270
rect 202 265 204 270
rect 196 254 198 257
rect 248 259 250 266
rect 202 254 204 255
rect 220 254 222 255
rect 229 254 231 257
rect 164 238 166 250
rect 170 247 172 250
rect 164 225 166 228
rect 248 252 250 255
rect 295 248 297 268
rect 305 248 307 268
rect 506 308 508 311
rect 683 327 685 330
rect 596 295 598 307
rect 636 301 638 313
rect 840 367 842 375
rect 778 348 780 351
rect 794 346 796 351
rect 788 335 790 338
rect 840 340 842 347
rect 794 335 796 336
rect 812 335 814 336
rect 821 335 823 338
rect 756 319 758 331
rect 762 328 764 331
rect 472 291 474 294
rect 482 291 484 294
rect 596 282 598 285
rect 393 279 395 282
rect 683 295 685 307
rect 723 301 725 313
rect 756 306 758 309
rect 683 282 685 285
rect 840 333 842 336
rect 840 320 842 323
rect 812 312 814 315
rect 821 312 823 315
rect 788 294 790 295
rect 794 292 796 295
rect 636 278 638 281
rect 723 278 725 281
rect 478 268 480 271
rect 488 268 490 271
rect 248 239 250 242
rect 220 231 222 234
rect 229 231 231 234
rect 358 241 360 259
rect 368 241 370 259
rect 393 245 395 259
rect 433 254 435 258
rect 443 254 445 258
rect 393 232 395 235
rect 358 228 360 231
rect 368 228 370 231
rect 295 224 297 228
rect 305 224 307 228
rect 433 215 435 234
rect 443 215 445 234
rect 690 254 692 257
rect 513 248 515 251
rect 756 252 758 255
rect 762 252 764 259
rect 778 252 780 264
rect 794 252 796 255
rect 196 213 198 214
rect 202 211 204 214
rect 358 201 360 204
rect 368 201 370 204
rect 46 179 48 182
rect 52 179 54 186
rect 68 179 70 191
rect 84 179 86 182
rect 130 175 132 183
rect 68 156 70 159
rect 84 154 86 159
rect 297 168 299 171
rect 307 168 309 171
rect 78 143 80 146
rect 130 148 132 155
rect 84 143 86 144
rect 102 143 104 144
rect 111 143 113 146
rect 46 127 48 139
rect 52 136 54 139
rect 46 114 48 117
rect 130 141 132 144
rect 130 128 132 131
rect 478 210 480 228
rect 488 210 490 228
rect 513 214 515 228
rect 690 222 692 234
rect 608 212 610 215
rect 840 248 842 256
rect 778 229 780 232
rect 794 227 796 232
rect 788 216 790 219
rect 840 221 842 228
rect 794 216 796 217
rect 812 216 814 217
rect 821 216 823 219
rect 513 201 515 204
rect 478 197 480 200
rect 488 197 490 200
rect 433 192 435 195
rect 443 192 445 195
rect 690 209 692 212
rect 705 203 707 204
rect 676 200 678 201
rect 608 180 610 192
rect 756 200 758 212
rect 762 209 764 212
rect 756 187 758 190
rect 705 180 707 183
rect 435 169 437 173
rect 445 169 447 173
rect 469 169 471 172
rect 676 177 678 180
rect 840 214 842 217
rect 840 201 842 204
rect 812 193 814 196
rect 821 193 823 196
rect 788 175 790 176
rect 720 170 722 173
rect 794 173 796 176
rect 358 143 360 161
rect 368 143 370 161
rect 608 167 610 170
rect 680 164 682 167
rect 623 161 625 162
rect 594 158 596 159
rect 358 130 360 133
rect 368 130 370 133
rect 435 130 437 149
rect 445 130 447 149
rect 469 137 471 149
rect 623 138 625 141
rect 102 120 104 123
rect 111 120 113 123
rect 297 109 299 128
rect 307 109 309 128
rect 352 111 354 114
rect 362 111 364 114
rect 78 102 80 103
rect 84 100 86 103
rect 161 92 163 95
rect 167 92 169 99
rect 183 92 185 104
rect 297 96 299 99
rect 307 96 309 99
rect 199 92 201 95
rect 245 88 247 96
rect 297 88 299 91
rect 307 88 309 91
rect 183 69 185 72
rect 199 67 201 72
rect 594 135 596 138
rect 680 132 682 144
rect 720 138 722 150
rect 638 128 640 131
rect 469 124 471 127
rect 598 122 600 125
rect 494 116 496 119
rect 504 116 506 119
rect 435 107 437 110
rect 445 107 447 110
rect 387 91 389 94
rect 411 90 413 94
rect 421 90 423 94
rect 193 56 195 59
rect 245 61 247 68
rect 199 56 201 57
rect 217 56 219 57
rect 226 56 228 59
rect 161 40 163 52
rect 167 49 169 52
rect 161 27 163 30
rect 245 54 247 57
rect 297 48 299 68
rect 307 48 309 68
rect 352 53 354 71
rect 362 53 364 71
rect 387 57 389 71
rect 680 119 682 122
rect 759 129 761 132
rect 765 129 767 136
rect 781 129 783 141
rect 797 129 799 132
rect 720 115 722 118
rect 529 96 531 99
rect 598 90 600 102
rect 638 96 640 108
rect 598 77 600 80
rect 843 125 845 133
rect 781 106 783 109
rect 797 104 799 109
rect 791 93 793 96
rect 843 98 845 105
rect 797 93 799 94
rect 815 93 817 94
rect 824 93 826 96
rect 759 77 761 89
rect 765 86 767 89
rect 245 41 247 44
rect 217 33 219 36
rect 226 33 228 36
rect 411 51 413 70
rect 421 51 423 70
rect 494 58 496 76
rect 504 58 506 76
rect 529 62 531 76
rect 638 73 640 76
rect 759 64 761 67
rect 387 44 389 47
rect 352 40 354 43
rect 362 40 364 43
rect 843 91 845 94
rect 843 78 845 81
rect 815 70 817 73
rect 824 70 826 73
rect 791 52 793 53
rect 529 49 531 52
rect 797 50 799 53
rect 494 45 496 48
rect 504 45 506 48
rect 411 28 413 31
rect 421 28 423 31
rect 297 24 299 28
rect 307 24 309 28
rect 193 15 195 16
rect 199 13 201 16
<< polycontact >>
rect 217 849 221 853
rect 265 839 269 843
rect 179 823 183 827
rect 496 832 500 836
rect 620 836 624 840
rect 668 826 672 830
rect 248 811 252 815
rect 484 810 488 814
rect 513 813 517 817
rect 213 793 217 797
rect 582 810 586 814
rect 651 798 655 802
rect 616 780 620 784
rect 217 738 221 742
rect 334 741 338 745
rect 344 734 348 738
rect 486 742 490 746
rect 265 728 269 732
rect 179 712 183 716
rect 104 678 108 682
rect 248 700 252 704
rect 213 682 217 686
rect 599 724 603 728
rect 678 730 682 734
rect 375 709 379 713
rect 587 702 591 706
rect 616 705 620 709
rect 666 708 670 712
rect 695 711 699 715
rect 152 668 156 672
rect 66 652 70 656
rect 297 657 301 661
rect 307 664 311 668
rect 135 640 139 644
rect 778 681 782 685
rect 826 671 830 675
rect 100 622 104 626
rect 207 599 211 603
rect 366 621 370 625
rect 376 627 380 631
rect 401 625 405 629
rect 589 634 593 638
rect 668 640 672 644
rect 740 655 744 659
rect 297 602 301 606
rect 307 610 311 614
rect 809 643 813 647
rect 774 625 778 629
rect 432 602 436 606
rect 255 589 259 593
rect 169 573 173 577
rect 96 537 100 541
rect 442 595 446 599
rect 238 561 242 565
rect 203 543 207 547
rect 144 527 148 531
rect 58 511 62 515
rect 127 499 131 503
rect 597 552 601 556
rect 688 552 692 556
rect 366 523 370 527
rect 376 529 380 533
rect 585 530 589 534
rect 614 533 618 537
rect 424 517 428 521
rect 434 510 438 514
rect 458 517 462 521
rect 92 481 96 485
rect 292 483 296 487
rect 302 490 306 494
rect 205 438 209 442
rect 676 530 680 534
rect 705 533 709 537
rect 253 428 257 432
rect 292 428 296 432
rect 167 412 171 416
rect 81 384 85 388
rect 302 436 306 440
rect 356 433 360 437
rect 366 439 370 443
rect 391 437 395 441
rect 587 462 591 466
rect 790 503 794 507
rect 838 493 842 497
rect 678 462 682 466
rect 752 477 756 481
rect 821 465 825 469
rect 786 447 790 451
rect 479 428 483 432
rect 489 434 493 438
rect 514 432 518 436
rect 236 400 240 404
rect 429 415 433 419
rect 439 408 443 412
rect 201 382 205 386
rect 129 374 133 378
rect 43 358 47 362
rect 112 346 116 350
rect 77 328 81 332
rect 602 386 606 390
rect 689 386 693 390
rect 590 364 594 368
rect 619 367 623 371
rect 347 335 351 339
rect 357 341 361 345
rect 291 310 295 314
rect 301 317 305 321
rect 677 364 681 368
rect 706 367 710 371
rect 468 322 472 326
rect 478 315 482 319
rect 502 322 506 326
rect 198 265 202 269
rect 246 255 250 259
rect 291 255 295 259
rect 160 239 164 243
rect 301 263 305 267
rect 592 296 596 300
rect 790 346 794 350
rect 838 336 842 340
rect 752 320 756 324
rect 679 296 683 300
rect 821 308 825 312
rect 786 290 790 294
rect 229 227 233 231
rect 354 242 358 246
rect 364 248 368 252
rect 389 246 393 250
rect 429 223 433 227
rect 439 216 443 220
rect 194 209 198 213
rect 80 154 84 158
rect 128 144 132 148
rect 42 128 46 132
rect 474 211 478 215
rect 484 217 488 221
rect 509 215 513 219
rect 686 223 690 227
rect 790 227 794 231
rect 838 217 842 221
rect 674 201 678 205
rect 703 204 707 208
rect 604 181 608 185
rect 752 201 756 205
rect 821 189 825 193
rect 786 171 790 175
rect 354 144 358 148
rect 364 150 368 154
rect 592 159 596 163
rect 621 162 625 166
rect 431 138 435 142
rect 441 131 445 135
rect 465 138 469 142
rect 111 116 115 120
rect 293 110 297 114
rect 303 117 307 121
rect 76 98 80 102
rect 195 67 199 71
rect 676 133 680 137
rect 243 57 247 61
rect 157 41 161 45
rect 293 55 297 59
rect 303 63 307 67
rect 348 54 352 58
rect 358 60 362 64
rect 383 58 387 62
rect 594 91 598 95
rect 793 104 797 108
rect 841 94 845 98
rect 755 78 759 82
rect 407 59 411 63
rect 226 29 230 33
rect 417 52 421 56
rect 490 59 494 63
rect 500 65 504 69
rect 525 63 529 67
rect 824 66 828 70
rect 789 48 793 52
rect 191 11 195 15
<< polynpluscontact >>
rect 526 748 530 752
rect 629 640 633 644
rect 708 646 712 650
rect 627 468 631 472
rect 718 468 722 472
rect 632 302 636 306
rect 719 302 723 306
rect 716 139 720 143
rect 634 97 638 101
<< metal1 >>
rect 15 898 327 901
rect 15 897 102 898
rect 15 606 19 897
rect 99 781 102 897
rect 200 892 203 898
rect 332 898 871 901
rect 178 889 265 892
rect 178 874 182 889
rect 200 874 204 889
rect 216 874 220 889
rect 262 870 265 889
rect 228 857 237 858
rect 228 854 261 857
rect 208 853 212 854
rect 208 849 217 853
rect 208 846 212 849
rect 204 843 214 846
rect 168 823 179 827
rect 192 825 196 834
rect 186 822 196 825
rect 178 792 182 812
rect 193 796 196 822
rect 204 815 207 843
rect 210 838 214 843
rect 232 838 235 854
rect 258 843 261 854
rect 272 843 276 850
rect 258 840 265 843
rect 272 839 322 843
rect 272 836 276 839
rect 204 811 248 815
rect 193 793 213 796
rect 181 790 182 792
rect 224 790 228 798
rect 255 790 258 818
rect 262 790 265 826
rect 181 787 265 790
rect 99 778 265 781
rect 99 777 182 778
rect 99 721 102 777
rect 178 763 182 777
rect 200 763 204 778
rect 216 763 220 778
rect 262 759 265 778
rect 228 746 237 747
rect 318 746 322 839
rect 342 782 345 898
rect 510 873 513 898
rect 590 879 593 898
rect 581 876 668 879
rect 474 870 528 873
rect 474 783 477 870
rect 495 863 498 870
rect 485 832 496 835
rect 504 835 507 843
rect 504 832 516 835
rect 480 814 483 832
rect 504 831 507 832
rect 495 817 498 821
rect 513 817 516 832
rect 495 814 500 817
rect 480 811 484 814
rect 519 789 522 792
rect 490 786 522 789
rect 333 779 372 782
rect 474 780 490 783
rect 333 772 336 779
rect 352 772 355 779
rect 228 743 261 746
rect 208 742 212 743
rect 208 738 217 742
rect 208 735 212 738
rect 204 732 214 735
rect 65 718 152 721
rect 65 703 69 718
rect 87 703 91 718
rect 103 703 107 718
rect 149 699 152 718
rect 167 712 179 716
rect 192 714 196 723
rect 186 711 196 714
rect 115 686 124 687
rect 115 683 148 686
rect 95 682 99 683
rect 95 678 104 682
rect 95 675 99 678
rect 91 672 101 675
rect 55 652 66 656
rect 79 654 83 663
rect 73 651 83 654
rect 65 621 69 641
rect 80 625 83 651
rect 91 644 94 672
rect 97 667 101 672
rect 119 667 122 683
rect 145 672 148 683
rect 159 672 163 679
rect 178 679 182 701
rect 193 685 196 711
rect 204 704 207 732
rect 210 727 214 732
rect 232 727 235 743
rect 258 732 261 743
rect 322 741 334 744
rect 343 744 346 752
rect 369 750 372 779
rect 485 773 488 780
rect 369 747 379 750
rect 343 741 361 744
rect 272 732 276 739
rect 305 733 315 737
rect 305 732 309 733
rect 320 734 344 737
rect 352 733 355 741
rect 258 729 265 732
rect 272 728 309 732
rect 272 725 276 728
rect 290 721 319 725
rect 296 715 300 721
rect 204 700 248 704
rect 193 682 213 685
rect 224 679 228 687
rect 255 679 258 707
rect 262 679 265 715
rect 333 710 336 713
rect 358 712 361 741
rect 374 740 377 747
rect 479 742 486 745
rect 494 745 497 753
rect 519 751 522 786
rect 525 779 528 870
rect 581 861 585 876
rect 603 861 607 876
rect 619 861 623 876
rect 665 857 668 876
rect 631 844 640 845
rect 631 841 664 844
rect 611 840 615 841
rect 611 836 620 840
rect 611 833 615 836
rect 607 830 617 833
rect 578 813 582 814
rect 562 810 582 813
rect 595 812 599 821
rect 519 748 526 751
rect 534 751 537 759
rect 562 751 565 810
rect 589 809 599 812
rect 581 777 585 799
rect 596 783 599 809
rect 607 802 610 830
rect 613 825 617 830
rect 635 825 638 841
rect 661 830 664 841
rect 675 830 679 837
rect 661 827 668 830
rect 675 826 691 830
rect 675 823 679 826
rect 607 798 651 802
rect 596 780 616 783
rect 627 777 631 785
rect 658 777 661 805
rect 665 779 668 813
rect 581 774 664 777
rect 707 771 710 898
rect 656 768 710 771
rect 656 765 659 768
rect 534 748 565 751
rect 577 762 659 765
rect 534 747 537 748
rect 494 742 509 745
rect 494 741 497 742
rect 485 724 488 731
rect 525 724 528 727
rect 485 721 500 724
rect 383 713 386 720
rect 505 721 528 724
rect 354 709 375 712
rect 383 710 423 713
rect 178 676 265 679
rect 145 669 152 672
rect 159 669 173 672
rect 159 668 165 669
rect 159 665 163 668
rect 91 640 135 644
rect 80 622 100 625
rect 111 619 115 627
rect 142 619 145 647
rect 149 649 152 655
rect 221 649 224 676
rect 149 646 224 649
rect 281 664 307 668
rect 149 619 152 646
rect 168 639 255 642
rect 281 640 284 664
rect 314 661 318 675
rect 168 635 172 639
rect 70 616 152 619
rect 158 631 172 635
rect 158 606 162 631
rect 168 624 172 631
rect 190 624 194 639
rect 206 624 210 639
rect 252 620 255 639
rect 15 602 162 606
rect 218 607 227 608
rect 218 604 251 607
rect 281 606 284 635
rect 287 657 297 661
rect 305 657 345 661
rect 305 656 309 657
rect 287 614 290 652
rect 296 642 300 646
rect 314 643 318 646
rect 314 642 330 643
rect 296 639 330 642
rect 296 635 300 639
rect 341 624 345 657
rect 358 631 361 709
rect 383 708 386 710
rect 374 694 377 698
rect 374 691 403 694
rect 510 694 513 721
rect 408 691 513 694
rect 365 685 398 688
rect 365 678 368 685
rect 395 668 398 685
rect 577 675 580 762
rect 598 755 601 762
rect 588 724 599 727
rect 607 727 610 735
rect 607 724 619 727
rect 583 706 586 724
rect 607 723 610 724
rect 598 709 601 713
rect 616 709 619 724
rect 598 706 603 709
rect 583 703 587 706
rect 622 681 625 684
rect 593 678 625 681
rect 577 672 593 675
rect 395 665 503 668
rect 400 658 403 665
rect 431 643 434 665
rect 358 628 376 631
rect 384 629 387 638
rect 409 629 412 638
rect 431 640 453 643
rect 431 633 434 640
rect 450 633 453 640
rect 384 626 401 629
rect 341 621 351 624
rect 356 621 366 624
rect 384 624 387 626
rect 409 626 418 629
rect 409 624 412 626
rect 374 621 387 624
rect 374 620 378 621
rect 287 610 307 614
rect 314 606 318 615
rect 198 603 202 604
rect 15 580 19 602
rect 198 599 207 603
rect 198 596 202 599
rect 194 593 204 596
rect 15 577 144 580
rect 15 576 61 577
rect 15 469 19 576
rect 57 562 61 576
rect 79 562 83 577
rect 95 562 99 577
rect 141 558 144 577
rect 155 573 169 577
rect 182 575 186 584
rect 176 572 186 575
rect 107 545 116 546
rect 107 542 140 545
rect 87 541 91 542
rect 87 537 96 541
rect 87 534 91 537
rect 83 531 93 534
rect 54 514 58 515
rect 47 511 58 514
rect 71 513 75 522
rect 65 510 75 513
rect 57 480 61 500
rect 72 484 75 510
rect 83 503 86 531
rect 89 526 93 531
rect 111 526 114 542
rect 137 531 140 542
rect 151 531 155 538
rect 168 540 172 562
rect 183 546 186 572
rect 194 565 197 593
rect 200 588 204 593
rect 222 588 225 604
rect 248 593 251 604
rect 262 593 266 600
rect 281 602 297 606
rect 305 602 340 606
rect 281 593 284 602
rect 248 590 255 593
rect 262 589 284 593
rect 305 595 309 602
rect 336 598 340 602
rect 365 604 368 610
rect 384 604 387 610
rect 400 606 403 614
rect 365 601 398 604
rect 415 605 418 626
rect 415 602 432 605
rect 441 605 444 613
rect 441 602 462 605
rect 333 595 442 598
rect 450 594 453 602
rect 363 589 398 592
rect 500 593 503 665
rect 588 665 591 672
rect 582 634 589 637
rect 597 637 600 645
rect 622 643 625 678
rect 628 671 631 762
rect 656 681 659 762
rect 677 761 680 768
rect 662 730 678 733
rect 686 733 689 741
rect 686 730 698 733
rect 662 721 665 730
rect 686 729 689 730
rect 662 712 665 716
rect 677 715 680 719
rect 695 715 698 730
rect 707 724 710 768
rect 760 727 765 732
rect 760 724 763 727
rect 707 721 826 724
rect 707 720 743 721
rect 677 712 682 715
rect 662 709 666 712
rect 701 687 704 690
rect 672 684 704 687
rect 656 678 672 681
rect 667 671 670 678
rect 622 640 629 643
rect 637 643 640 651
rect 637 640 656 643
rect 637 639 640 640
rect 597 634 612 637
rect 661 640 668 643
rect 676 643 679 651
rect 701 649 704 684
rect 707 677 710 720
rect 739 706 743 720
rect 760 716 765 721
rect 761 706 765 716
rect 777 706 781 721
rect 823 702 826 721
rect 789 689 798 690
rect 789 686 822 689
rect 769 685 773 686
rect 769 681 778 685
rect 769 678 773 681
rect 765 675 775 678
rect 701 646 708 649
rect 716 649 719 657
rect 732 655 740 659
rect 753 657 757 666
rect 732 649 735 655
rect 747 654 757 657
rect 716 646 735 649
rect 716 645 719 646
rect 676 640 691 643
rect 676 639 679 640
rect 597 633 600 634
rect 588 616 591 623
rect 667 622 670 629
rect 707 622 710 625
rect 739 622 743 644
rect 754 628 757 654
rect 765 647 768 675
rect 771 670 775 675
rect 793 670 796 686
rect 819 675 822 686
rect 833 675 837 682
rect 819 672 826 675
rect 833 671 847 675
rect 833 668 837 671
rect 765 643 809 647
rect 754 625 774 628
rect 785 622 789 630
rect 816 622 819 650
rect 823 624 826 658
rect 667 619 682 622
rect 628 616 631 619
rect 667 616 670 619
rect 687 619 822 622
rect 591 613 603 616
rect 608 613 670 616
rect 868 593 871 898
rect 498 590 871 593
rect 262 586 266 589
rect 365 580 368 589
rect 395 586 398 589
rect 498 586 501 590
rect 395 583 501 586
rect 194 561 238 565
rect 183 543 203 546
rect 214 540 218 548
rect 245 540 248 568
rect 252 540 255 576
rect 296 567 300 575
rect 314 569 318 575
rect 314 567 319 569
rect 296 564 319 567
rect 395 558 398 583
rect 417 574 431 578
rect 431 568 434 574
rect 395 555 460 558
rect 168 537 255 540
rect 266 548 314 551
rect 137 528 144 531
rect 151 530 157 531
rect 151 527 170 530
rect 151 524 155 527
rect 83 499 127 503
rect 72 481 92 484
rect 103 478 107 486
rect 134 478 137 506
rect 141 497 144 514
rect 214 497 217 537
rect 141 494 217 497
rect 141 478 144 494
rect 266 481 269 548
rect 285 547 314 548
rect 423 548 426 555
rect 442 548 445 555
rect 291 541 295 547
rect 457 548 460 555
rect 357 530 376 533
rect 384 531 387 540
rect 384 528 395 531
rect 321 523 337 526
rect 342 523 366 526
rect 384 526 387 528
rect 374 523 387 526
rect 61 475 144 478
rect 166 478 269 481
rect 276 490 302 494
rect 166 469 170 478
rect 15 465 170 469
rect 15 427 19 465
rect 166 463 170 465
rect 188 463 192 478
rect 204 463 208 478
rect 250 459 253 478
rect 276 467 279 490
rect 309 487 313 501
rect 321 487 324 523
rect 216 446 225 447
rect 216 443 249 446
rect 196 442 200 443
rect 196 438 205 442
rect 196 435 200 438
rect 192 432 202 435
rect 15 424 129 427
rect 15 423 46 424
rect 15 308 19 423
rect 42 409 46 423
rect 64 409 68 424
rect 80 409 84 424
rect 126 405 129 424
rect 151 412 167 416
rect 180 414 184 423
rect 174 411 184 414
rect 92 392 101 393
rect 92 389 125 392
rect 72 388 76 389
rect 72 384 81 388
rect 72 381 76 384
rect 68 378 78 381
rect 31 358 43 362
rect 56 360 60 369
rect 50 357 60 360
rect 42 327 46 347
rect 57 331 60 357
rect 68 350 71 378
rect 74 373 78 378
rect 96 373 99 389
rect 122 378 125 389
rect 136 378 140 385
rect 166 379 170 401
rect 181 385 184 411
rect 192 404 195 432
rect 198 427 202 432
rect 220 427 223 443
rect 246 432 249 443
rect 260 432 264 439
rect 276 432 279 462
rect 287 483 292 487
rect 300 483 324 487
rect 300 482 304 483
rect 282 440 285 482
rect 291 468 295 472
rect 309 468 313 472
rect 291 465 313 468
rect 291 461 295 465
rect 300 454 303 465
rect 282 436 302 440
rect 309 432 313 441
rect 348 443 351 523
rect 374 522 378 523
rect 365 508 368 512
rect 366 506 368 508
rect 384 506 387 512
rect 392 513 395 528
rect 413 517 424 520
rect 433 520 436 528
rect 466 521 469 528
rect 433 517 458 520
rect 466 518 475 521
rect 392 510 434 513
rect 442 509 445 517
rect 466 516 469 518
rect 366 503 411 506
rect 355 497 388 500
rect 355 490 358 497
rect 385 480 388 497
rect 408 486 411 503
rect 423 486 426 489
rect 457 486 460 506
rect 408 483 460 486
rect 385 477 431 480
rect 390 470 393 477
rect 428 456 431 477
rect 348 440 366 443
rect 374 441 377 450
rect 399 441 402 450
rect 428 453 450 456
rect 428 446 431 453
rect 447 446 450 453
rect 374 438 391 441
rect 335 433 356 436
rect 374 436 377 438
rect 399 438 408 441
rect 472 438 475 518
rect 498 509 501 583
rect 498 495 501 504
rect 575 503 578 590
rect 596 583 599 590
rect 586 552 597 555
rect 605 555 608 563
rect 605 552 617 555
rect 581 534 584 552
rect 605 551 608 552
rect 596 537 599 541
rect 614 537 617 552
rect 596 534 601 537
rect 581 531 585 534
rect 620 509 623 512
rect 591 506 623 509
rect 575 500 591 503
rect 478 492 511 495
rect 478 485 481 492
rect 508 475 511 492
rect 586 493 589 500
rect 508 472 516 475
rect 513 465 516 472
rect 580 462 587 465
rect 595 465 598 473
rect 620 471 623 506
rect 626 499 629 590
rect 666 503 669 590
rect 687 583 690 590
rect 677 552 688 555
rect 696 555 699 563
rect 696 552 708 555
rect 672 534 675 552
rect 696 551 699 552
rect 687 537 690 541
rect 705 537 708 552
rect 687 534 692 537
rect 672 531 676 534
rect 711 509 714 512
rect 682 506 714 509
rect 666 500 682 503
rect 677 493 680 500
rect 620 468 627 471
rect 635 471 638 479
rect 635 468 644 471
rect 635 467 638 468
rect 595 462 610 465
rect 641 465 644 468
rect 641 462 666 465
rect 595 461 598 462
rect 671 462 678 465
rect 686 465 689 473
rect 711 471 714 506
rect 717 499 720 590
rect 868 546 871 590
rect 751 543 871 546
rect 751 528 755 543
rect 773 528 777 543
rect 789 528 793 543
rect 835 524 838 543
rect 801 511 810 512
rect 801 508 834 511
rect 781 507 785 508
rect 781 503 790 507
rect 781 500 785 503
rect 777 497 787 500
rect 711 468 718 471
rect 726 471 729 479
rect 742 477 752 481
rect 765 479 769 488
rect 742 471 745 477
rect 759 476 769 479
rect 726 468 745 471
rect 726 467 729 468
rect 686 462 701 465
rect 686 461 689 462
rect 399 436 402 438
rect 365 433 377 436
rect 365 432 368 433
rect 246 429 253 432
rect 260 428 292 432
rect 300 428 325 432
rect 260 425 264 428
rect 300 421 304 428
rect 192 400 236 404
rect 181 382 201 385
rect 212 379 216 387
rect 243 379 246 407
rect 250 379 253 415
rect 322 410 325 428
rect 355 421 358 422
rect 353 416 358 421
rect 374 416 377 422
rect 390 418 393 426
rect 405 418 408 438
rect 471 435 489 438
rect 497 436 500 445
rect 522 436 525 445
rect 586 444 589 451
rect 626 444 629 447
rect 677 444 680 451
rect 717 444 720 447
rect 751 444 755 466
rect 766 450 769 476
rect 777 469 780 497
rect 783 492 787 497
rect 805 492 808 508
rect 831 497 834 508
rect 845 497 849 504
rect 831 494 838 497
rect 845 493 858 497
rect 845 490 849 493
rect 777 465 821 469
rect 766 447 786 450
rect 797 444 801 452
rect 828 444 831 472
rect 835 446 838 480
rect 586 441 601 444
rect 606 441 692 444
rect 697 441 834 444
rect 497 433 514 436
rect 355 413 390 416
rect 405 415 429 418
rect 438 418 441 426
rect 467 428 479 431
rect 497 431 500 433
rect 522 433 531 436
rect 522 431 525 433
rect 488 428 500 431
rect 467 418 470 428
rect 488 427 491 428
rect 868 427 871 543
rect 580 424 871 427
rect 438 415 470 418
rect 322 407 346 410
rect 421 410 439 411
rect 351 408 439 410
rect 351 407 424 408
rect 447 407 450 415
rect 291 393 295 401
rect 344 401 387 404
rect 478 411 481 417
rect 497 411 500 417
rect 513 413 516 421
rect 478 408 513 411
rect 309 395 313 401
rect 309 393 314 395
rect 291 390 314 393
rect 346 392 349 401
rect 122 375 129 378
rect 136 377 142 378
rect 136 374 154 377
rect 166 376 253 379
rect 136 371 140 374
rect 68 346 112 350
rect 57 328 77 331
rect 88 325 92 333
rect 119 325 122 353
rect 126 326 129 361
rect 203 326 206 376
rect 284 374 313 378
rect 290 371 294 374
rect 126 325 206 326
rect 47 323 206 325
rect 243 368 294 371
rect 47 322 129 323
rect 243 308 246 368
rect 384 363 387 401
rect 428 384 431 387
rect 478 384 481 408
rect 428 381 481 384
rect 580 363 583 424
rect 601 417 604 424
rect 591 386 602 389
rect 610 389 613 397
rect 610 386 622 389
rect 586 368 589 386
rect 610 385 613 386
rect 601 371 604 375
rect 619 371 622 386
rect 601 368 606 371
rect 586 365 590 368
rect 384 360 583 363
rect 338 342 357 345
rect 365 343 368 352
rect 384 351 387 360
rect 467 353 470 360
rect 486 353 489 360
rect 501 353 504 360
rect 365 340 418 343
rect 321 335 347 338
rect 365 338 368 340
rect 356 335 368 338
rect 15 305 246 308
rect 15 304 163 305
rect 15 197 19 304
rect 159 290 163 304
rect 181 290 185 305
rect 197 290 201 305
rect 243 286 246 305
rect 275 317 301 321
rect 275 301 278 317
rect 308 314 312 328
rect 321 314 325 335
rect 209 273 218 274
rect 209 270 242 273
rect 189 269 193 270
rect 189 265 198 269
rect 189 262 193 265
rect 185 259 195 262
rect 143 239 160 243
rect 173 241 177 250
rect 167 238 177 241
rect 159 208 163 228
rect 174 212 177 238
rect 185 231 188 259
rect 191 254 195 259
rect 213 254 216 270
rect 239 259 242 270
rect 253 259 257 266
rect 275 259 278 296
rect 286 310 291 314
rect 299 310 325 314
rect 299 309 303 310
rect 281 267 284 309
rect 290 295 294 299
rect 308 295 312 299
rect 290 292 312 295
rect 290 288 294 292
rect 299 281 302 292
rect 281 263 301 267
rect 308 259 312 268
rect 239 256 246 259
rect 253 255 291 259
rect 299 255 322 259
rect 253 252 257 255
rect 299 248 303 255
rect 334 245 337 335
rect 356 334 359 335
rect 346 318 349 324
rect 365 318 368 324
rect 346 315 373 318
rect 383 309 386 331
rect 415 318 418 340
rect 580 337 583 360
rect 625 343 628 346
rect 596 340 628 343
rect 580 334 596 337
rect 459 322 468 325
rect 477 325 480 333
rect 510 326 513 333
rect 591 327 594 334
rect 477 322 502 325
rect 510 323 519 326
rect 415 315 478 318
rect 486 314 489 322
rect 510 321 513 323
rect 353 306 386 309
rect 353 299 356 306
rect 383 289 386 306
rect 383 286 432 289
rect 467 291 470 294
rect 501 291 504 311
rect 462 288 504 291
rect 388 279 391 286
rect 428 264 432 286
rect 516 285 519 323
rect 585 296 592 299
rect 600 299 603 307
rect 625 305 628 340
rect 631 333 634 424
rect 667 337 670 424
rect 688 417 691 424
rect 678 386 689 389
rect 697 389 700 397
rect 697 386 709 389
rect 673 368 676 386
rect 697 385 700 386
rect 688 371 691 375
rect 706 371 709 386
rect 688 368 693 371
rect 673 365 677 368
rect 712 343 715 346
rect 683 340 715 343
rect 667 334 683 337
rect 678 327 681 334
rect 625 302 632 305
rect 640 305 643 313
rect 640 302 662 305
rect 640 301 643 302
rect 600 296 615 299
rect 659 299 662 302
rect 659 296 667 299
rect 600 295 603 296
rect 672 296 679 299
rect 687 299 690 307
rect 712 305 715 340
rect 718 333 721 424
rect 868 389 871 424
rect 751 386 871 389
rect 751 371 755 386
rect 773 371 777 386
rect 789 371 793 386
rect 835 367 838 386
rect 801 354 810 355
rect 801 351 834 354
rect 781 350 785 351
rect 781 346 790 350
rect 781 343 785 346
rect 777 340 787 343
rect 744 320 752 324
rect 765 322 769 331
rect 712 302 719 305
rect 727 305 730 313
rect 744 305 747 320
rect 759 319 769 322
rect 727 302 747 305
rect 727 301 730 302
rect 687 296 702 299
rect 687 295 690 296
rect 467 282 519 285
rect 751 287 755 309
rect 766 293 769 319
rect 777 312 780 340
rect 783 335 787 340
rect 805 335 808 351
rect 831 340 834 351
rect 845 340 849 347
rect 831 337 838 340
rect 845 336 860 340
rect 845 333 849 336
rect 777 308 821 312
rect 766 290 786 293
rect 797 287 801 295
rect 828 287 831 315
rect 835 289 838 323
rect 345 249 364 252
rect 372 250 375 259
rect 397 250 400 259
rect 428 261 450 264
rect 428 254 431 261
rect 447 254 450 261
rect 372 247 389 250
rect 334 242 354 245
rect 372 245 375 247
rect 397 247 406 250
rect 397 245 400 247
rect 363 242 375 245
rect 185 227 229 231
rect 174 209 194 212
rect 205 206 209 214
rect 236 206 239 234
rect 243 206 246 242
rect 290 220 294 228
rect 308 222 312 228
rect 308 220 313 222
rect 290 217 313 220
rect 164 203 246 206
rect 15 194 128 197
rect 15 193 45 194
rect 15 84 19 193
rect 41 179 45 193
rect 63 179 67 194
rect 79 179 83 194
rect 125 189 128 194
rect 125 186 289 189
rect 125 175 128 186
rect 286 178 289 186
rect 286 174 315 178
rect 292 168 296 174
rect 91 162 100 163
rect 91 159 124 162
rect 71 158 75 159
rect 71 154 80 158
rect 71 151 75 154
rect 67 148 77 151
rect 25 128 42 132
rect 55 130 59 139
rect 49 127 59 130
rect 41 97 45 117
rect 56 101 59 127
rect 67 120 70 148
rect 73 143 77 148
rect 95 143 98 159
rect 121 148 124 159
rect 135 148 139 155
rect 334 154 337 242
rect 363 241 366 242
rect 353 225 356 231
rect 372 225 375 231
rect 388 225 391 235
rect 353 222 394 225
rect 403 226 406 247
rect 403 223 429 226
rect 438 226 441 234
rect 438 223 456 226
rect 346 216 439 219
rect 447 215 450 223
rect 351 210 390 213
rect 453 214 456 223
rect 467 221 470 282
rect 591 278 594 285
rect 631 278 634 281
rect 678 278 681 285
rect 751 284 834 287
rect 718 278 721 281
rect 751 278 754 284
rect 473 275 506 278
rect 591 275 606 278
rect 473 268 476 275
rect 503 258 506 275
rect 611 275 693 278
rect 698 275 754 278
rect 751 269 838 270
rect 868 269 871 386
rect 751 267 871 269
rect 751 264 755 267
rect 618 261 755 264
rect 618 258 621 261
rect 503 255 621 258
rect 508 248 511 255
rect 467 218 484 221
rect 492 219 495 228
rect 517 219 520 228
rect 618 222 621 255
rect 492 216 509 219
rect 453 211 474 214
rect 492 214 495 216
rect 517 216 524 219
rect 582 219 636 222
rect 517 214 520 216
rect 483 211 495 214
rect 483 210 486 211
rect 353 201 356 210
rect 387 176 390 210
rect 428 192 431 195
rect 473 194 476 200
rect 492 194 495 200
rect 508 194 511 204
rect 466 192 543 194
rect 425 191 543 192
rect 425 189 469 191
rect 582 179 585 219
rect 603 212 606 219
rect 395 176 585 179
rect 430 169 433 176
rect 449 169 452 176
rect 464 169 467 176
rect 334 151 364 154
rect 372 152 375 161
rect 372 149 407 152
rect 121 145 128 148
rect 135 144 150 148
rect 334 144 354 147
rect 372 147 375 149
rect 363 144 375 147
rect 135 141 139 144
rect 67 116 111 120
rect 56 98 76 101
rect 87 95 91 103
rect 118 95 121 123
rect 125 95 128 131
rect 277 117 303 121
rect 156 107 243 110
rect 156 105 160 107
rect 46 92 128 95
rect 140 101 160 105
rect 140 84 144 101
rect 156 92 160 101
rect 178 92 182 107
rect 194 92 198 107
rect 240 88 243 107
rect 277 96 280 117
rect 310 114 314 128
rect 334 114 337 144
rect 363 143 366 144
rect 353 127 356 133
rect 372 127 375 133
rect 404 134 407 149
rect 423 138 431 141
rect 440 141 443 149
rect 473 142 476 149
rect 440 138 465 141
rect 473 139 482 142
rect 404 131 441 134
rect 449 130 452 138
rect 473 137 476 139
rect 353 124 407 127
rect 15 80 144 84
rect 206 75 215 76
rect 206 72 239 75
rect 186 71 190 72
rect 186 67 195 71
rect 186 64 190 67
rect 182 61 192 64
rect 137 41 157 45
rect 170 43 174 52
rect 164 40 174 43
rect 156 8 160 30
rect 171 14 174 40
rect 182 33 185 61
rect 188 56 192 61
rect 210 56 213 72
rect 236 61 239 72
rect 250 61 254 68
rect 277 61 280 91
rect 288 110 293 114
rect 301 110 337 114
rect 301 109 305 110
rect 283 67 286 109
rect 292 95 296 99
rect 310 95 314 99
rect 292 92 314 95
rect 292 88 296 92
rect 301 83 304 92
rect 334 80 337 110
rect 347 118 380 121
rect 347 111 350 118
rect 377 101 380 118
rect 404 107 407 124
rect 430 107 433 110
rect 464 107 467 127
rect 404 104 452 107
rect 457 104 467 107
rect 377 100 385 101
rect 377 98 390 100
rect 382 97 390 98
rect 395 97 428 100
rect 382 91 385 97
rect 406 90 409 97
rect 425 90 428 97
rect 326 77 337 80
rect 283 63 303 67
rect 236 58 243 61
rect 250 59 280 61
rect 310 59 314 68
rect 250 57 293 59
rect 250 54 254 57
rect 277 55 293 57
rect 301 55 320 59
rect 301 48 305 55
rect 182 29 226 33
rect 171 11 191 14
rect 202 8 206 16
rect 233 8 236 36
rect 240 10 243 44
rect 292 20 296 28
rect 310 22 314 28
rect 317 28 320 55
rect 326 57 329 77
rect 338 61 358 64
rect 366 62 369 71
rect 391 62 394 71
rect 366 59 383 62
rect 326 54 348 57
rect 366 57 369 59
rect 391 59 407 62
rect 416 62 419 70
rect 479 69 482 139
rect 489 126 492 176
rect 582 132 585 176
rect 593 181 604 184
rect 612 184 615 192
rect 612 181 624 184
rect 612 180 615 181
rect 588 163 591 179
rect 603 166 606 170
rect 621 166 624 181
rect 633 174 636 219
rect 664 185 667 261
rect 685 254 688 261
rect 670 223 686 226
rect 694 226 697 234
rect 694 223 706 226
rect 670 220 673 223
rect 694 222 697 223
rect 670 205 673 215
rect 685 208 688 212
rect 703 208 706 223
rect 685 205 690 208
rect 670 202 674 205
rect 709 180 712 183
rect 680 177 712 180
rect 633 171 680 174
rect 603 163 608 166
rect 588 160 592 163
rect 627 138 630 141
rect 598 135 630 138
rect 582 129 598 132
rect 489 123 522 126
rect 489 116 492 123
rect 519 106 522 123
rect 593 122 596 129
rect 519 103 527 106
rect 524 96 527 103
rect 587 91 594 94
rect 602 94 605 102
rect 627 100 630 135
rect 633 128 636 171
rect 675 164 678 171
rect 669 133 676 136
rect 684 136 687 144
rect 709 142 712 177
rect 715 170 718 261
rect 751 252 755 261
rect 773 252 777 267
rect 789 252 793 267
rect 835 266 871 267
rect 835 248 838 266
rect 801 235 810 236
rect 801 232 834 235
rect 781 231 785 232
rect 781 227 790 231
rect 781 224 785 227
rect 777 221 787 224
rect 742 202 752 205
rect 709 139 716 142
rect 724 142 727 150
rect 742 142 745 202
rect 748 201 752 202
rect 765 203 769 212
rect 759 200 769 203
rect 751 168 755 190
rect 766 174 769 200
rect 777 193 780 221
rect 783 216 787 221
rect 805 216 808 232
rect 831 221 834 232
rect 845 221 849 228
rect 831 218 838 221
rect 845 217 862 221
rect 845 214 849 217
rect 777 189 821 193
rect 766 171 786 174
rect 797 168 801 176
rect 828 168 831 196
rect 835 170 838 204
rect 751 165 834 168
rect 868 147 871 266
rect 724 139 745 142
rect 754 144 871 147
rect 724 138 727 139
rect 684 133 699 136
rect 684 132 687 133
rect 627 97 634 100
rect 642 100 645 108
rect 664 100 667 131
rect 754 129 758 144
rect 776 129 780 144
rect 792 129 796 144
rect 838 125 841 144
rect 675 115 678 122
rect 715 115 718 118
rect 675 112 690 115
rect 695 112 718 115
rect 804 112 813 113
rect 804 109 837 112
rect 784 108 788 109
rect 784 104 793 108
rect 784 101 788 104
rect 642 97 667 100
rect 780 98 790 101
rect 642 96 645 97
rect 602 91 617 94
rect 602 90 605 91
rect 479 66 500 69
rect 508 67 511 76
rect 533 67 536 76
rect 593 73 596 80
rect 746 78 755 82
rect 768 80 772 89
rect 633 73 636 76
rect 593 70 608 73
rect 613 70 636 73
rect 508 64 525 67
rect 416 59 490 62
rect 508 62 511 64
rect 533 64 544 67
rect 533 62 536 64
rect 499 59 511 62
rect 391 57 394 59
rect 357 54 369 57
rect 357 53 360 54
rect 397 52 417 55
rect 347 37 350 43
rect 366 37 369 43
rect 347 34 373 37
rect 382 37 385 47
rect 378 34 385 37
rect 397 28 400 52
rect 425 51 428 59
rect 499 58 502 59
rect 541 60 544 64
rect 746 60 749 78
rect 762 77 772 80
rect 541 57 749 60
rect 489 42 492 48
rect 508 42 511 48
rect 489 39 514 42
rect 524 42 527 52
rect 754 45 758 67
rect 769 51 772 77
rect 780 70 783 98
rect 786 93 790 98
rect 808 93 811 109
rect 834 98 837 109
rect 848 98 852 105
rect 834 95 841 98
rect 848 94 867 98
rect 848 91 852 94
rect 780 66 824 70
rect 769 48 789 51
rect 800 45 804 53
rect 831 45 834 73
rect 838 47 841 81
rect 754 42 837 45
rect 519 39 527 42
rect 406 28 409 31
rect 317 25 400 28
rect 310 20 315 22
rect 292 17 315 20
rect 156 5 240 8
<< m2contact >>
rect 327 896 332 901
rect 176 787 181 792
rect 500 812 505 817
rect 319 721 324 726
rect 664 774 669 779
rect 509 742 514 747
rect 500 719 505 724
rect 332 705 337 710
rect 423 710 428 715
rect 173 667 178 672
rect 65 616 70 621
rect 330 639 335 644
rect 403 691 408 696
rect 603 704 608 709
rect 351 619 356 624
rect 398 601 403 606
rect 462 602 467 607
rect 328 593 333 598
rect 662 716 667 721
rect 682 710 687 715
rect 612 634 617 639
rect 656 638 661 643
rect 691 640 696 645
rect 682 617 687 622
rect 822 619 827 624
rect 603 611 608 616
rect 319 564 324 569
rect 412 573 417 578
rect 170 525 175 530
rect 56 475 61 480
rect 314 547 319 552
rect 352 530 357 535
rect 337 523 342 528
rect 361 503 366 508
rect 330 433 335 438
rect 601 532 606 537
rect 672 552 677 557
rect 692 532 697 537
rect 610 462 615 467
rect 666 460 671 465
rect 701 462 706 467
rect 601 439 606 444
rect 692 439 697 444
rect 834 441 839 446
rect 390 413 395 418
rect 531 433 536 438
rect 346 407 351 412
rect 314 390 319 395
rect 151 369 156 374
rect 42 322 47 327
rect 313 374 318 379
rect 423 381 428 386
rect 606 366 611 371
rect 333 342 338 347
rect 383 346 388 351
rect 299 276 304 281
rect 322 255 327 260
rect 383 331 388 336
rect 373 315 378 320
rect 454 322 459 327
rect 457 288 462 293
rect 673 386 678 391
rect 693 366 698 371
rect 615 296 620 301
rect 667 294 672 299
rect 702 296 707 301
rect 340 249 345 254
rect 159 203 164 208
rect 313 217 318 222
rect 315 174 320 179
rect 394 222 399 227
rect 340 216 346 222
rect 834 284 839 289
rect 606 273 611 278
rect 693 273 698 278
rect 420 189 425 194
rect 543 191 548 196
rect 390 174 395 179
rect 150 144 155 149
rect 41 92 46 97
rect 418 138 423 143
rect 301 78 306 83
rect 452 102 457 107
rect 390 97 395 102
rect 333 61 338 66
rect 690 203 695 208
rect 608 161 613 166
rect 664 131 669 136
rect 834 165 839 170
rect 699 133 704 138
rect 690 110 695 115
rect 617 91 622 96
rect 608 68 613 73
rect 373 34 378 39
rect 514 39 519 44
rect 837 42 842 47
rect 405 23 410 28
rect 315 17 320 22
rect 240 5 245 10
<< pm12contact >>
rect 189 881 194 886
rect 207 881 212 886
rect 221 839 226 844
rect 239 839 244 844
rect 189 770 194 775
rect 207 770 212 775
rect 76 710 81 715
rect 94 710 99 715
rect 108 668 113 673
rect 126 668 131 673
rect 221 728 226 733
rect 239 728 244 733
rect 592 868 597 873
rect 610 868 615 873
rect 624 826 629 831
rect 642 826 647 831
rect 179 631 184 636
rect 197 631 202 636
rect 68 569 73 574
rect 86 569 91 574
rect 100 527 105 532
rect 118 527 123 532
rect 211 589 216 594
rect 229 589 234 594
rect 750 713 755 718
rect 768 713 773 718
rect 782 671 787 676
rect 800 671 805 676
rect 177 470 182 475
rect 195 470 200 475
rect 53 416 58 421
rect 71 416 76 421
rect 85 374 90 379
rect 103 374 108 379
rect 209 428 214 433
rect 227 428 232 433
rect 762 535 767 540
rect 780 535 785 540
rect 794 493 799 498
rect 812 493 817 498
rect 170 297 175 302
rect 188 297 193 302
rect 202 255 207 260
rect 220 255 225 260
rect 762 378 767 383
rect 780 378 785 383
rect 794 336 799 341
rect 812 336 817 341
rect 52 186 57 191
rect 70 186 75 191
rect 84 144 89 149
rect 102 144 107 149
rect 167 99 172 104
rect 185 99 190 104
rect 199 57 204 62
rect 217 57 222 62
rect 762 259 767 264
rect 780 259 785 264
rect 794 217 799 222
rect 812 217 817 222
rect 765 136 770 141
rect 783 136 788 141
rect 797 94 802 99
rect 815 94 820 99
<< psm12contact >>
rect 408 517 413 522
<< ndm12contact >>
rect 480 789 485 794
rect 509 792 514 797
rect 583 681 588 686
rect 612 684 617 689
rect 662 687 667 692
rect 691 690 696 695
rect 581 509 586 514
rect 610 512 615 517
rect 672 509 677 514
rect 701 512 706 517
rect 586 343 591 348
rect 615 346 620 351
rect 673 343 678 348
rect 702 346 707 351
rect 670 180 675 185
rect 699 183 704 188
rect 588 138 593 143
rect 617 141 622 146
<< metal2 >>
rect 7 906 884 909
rect 78 881 189 884
rect 194 881 207 884
rect 7 790 10 879
rect 197 842 200 881
rect 197 839 221 842
rect 226 839 239 842
rect 7 787 176 790
rect 7 619 10 787
rect 77 770 189 773
rect 194 770 207 773
rect 197 731 200 770
rect 197 728 221 731
rect 226 728 239 731
rect 327 726 330 896
rect 324 723 330 726
rect 81 710 94 713
rect 84 671 87 710
rect 84 668 108 671
rect 113 668 126 671
rect 7 616 65 619
rect 7 478 10 616
rect 84 594 87 668
rect 175 657 178 667
rect 175 654 287 657
rect 184 631 197 634
rect 187 592 190 631
rect 89 589 211 592
rect 216 589 229 592
rect 73 569 86 572
rect 321 569 324 721
rect 332 696 335 705
rect 405 696 408 906
rect 602 871 605 886
rect 597 868 610 871
rect 600 829 603 868
rect 600 826 624 829
rect 629 826 642 829
rect 474 789 480 794
rect 474 745 477 789
rect 502 724 505 812
rect 509 747 512 792
rect 881 777 884 906
rect 669 774 884 777
rect 553 716 662 719
rect 332 693 403 696
rect 333 665 336 693
rect 553 713 556 716
rect 428 710 556 713
rect 760 716 763 727
rect 755 713 768 716
rect 330 662 336 665
rect 330 644 333 662
rect 76 530 79 569
rect 76 527 100 530
rect 105 527 118 530
rect 7 475 56 478
rect 7 325 10 475
rect 76 433 79 527
rect 172 486 175 525
rect 172 483 282 486
rect 182 470 195 473
rect 185 431 188 470
rect 81 428 209 431
rect 214 428 227 431
rect 58 416 71 419
rect 61 377 64 416
rect 316 395 319 547
rect 330 438 333 593
rect 353 535 356 619
rect 403 577 407 606
rect 403 573 412 577
rect 423 532 426 710
rect 577 681 583 686
rect 577 637 580 681
rect 605 616 608 704
rect 656 687 662 692
rect 612 639 615 684
rect 656 643 659 687
rect 684 622 687 710
rect 691 645 694 690
rect 758 674 761 713
rect 758 671 782 674
rect 787 671 800 674
rect 881 622 884 774
rect 827 619 884 622
rect 464 580 467 602
rect 464 577 675 580
rect 408 529 426 532
rect 61 374 85 377
rect 90 374 103 377
rect 7 322 42 325
rect 7 288 10 322
rect 7 206 10 283
rect 61 260 64 374
rect 151 313 154 369
rect 151 310 281 313
rect 175 297 188 300
rect 178 258 181 297
rect 267 276 299 279
rect 66 255 202 258
rect 207 255 220 258
rect 7 203 159 206
rect 7 3 10 203
rect 57 186 70 189
rect 60 147 63 186
rect 60 144 84 147
rect 89 144 102 147
rect 41 3 44 92
rect 60 62 63 144
rect 152 114 155 144
rect 267 128 270 276
rect 315 222 318 374
rect 339 352 342 523
rect 408 522 411 529
rect 348 505 361 508
rect 348 421 351 505
rect 333 349 342 352
rect 333 347 339 349
rect 348 257 351 407
rect 392 384 395 413
rect 392 381 423 384
rect 383 336 386 346
rect 464 334 467 577
rect 672 557 675 577
rect 771 538 774 551
rect 767 535 780 538
rect 575 509 581 514
rect 575 465 578 509
rect 603 444 606 532
rect 610 467 613 512
rect 666 509 672 514
rect 666 465 669 509
rect 694 444 697 532
rect 701 467 704 512
rect 770 496 773 535
rect 770 493 794 496
rect 799 493 812 496
rect 881 444 884 619
rect 839 441 884 444
rect 456 331 467 334
rect 533 404 536 433
rect 881 413 884 441
rect 533 401 676 404
rect 456 327 459 331
rect 378 315 403 318
rect 400 293 403 315
rect 400 290 457 293
rect 324 219 327 255
rect 340 254 351 257
rect 324 216 340 219
rect 152 111 283 114
rect 172 99 185 102
rect 175 60 178 99
rect 65 57 199 60
rect 204 57 217 60
rect 240 3 245 5
rect 301 3 304 78
rect 317 22 320 174
rect 340 76 343 216
rect 396 192 399 222
rect 396 189 420 192
rect 533 185 536 401
rect 673 391 676 401
rect 771 381 774 393
rect 767 378 780 381
rect 580 343 586 348
rect 580 299 583 343
rect 608 278 611 366
rect 615 301 618 346
rect 667 343 673 348
rect 667 299 670 343
rect 695 278 698 366
rect 702 301 705 346
rect 770 339 773 378
rect 770 336 794 339
rect 799 336 812 339
rect 881 287 884 408
rect 839 284 884 287
rect 771 262 774 274
rect 767 259 780 262
rect 770 220 773 259
rect 770 217 794 220
rect 799 217 812 220
rect 418 182 536 185
rect 390 102 393 174
rect 418 143 421 182
rect 335 73 343 76
rect 335 66 338 73
rect 375 3 378 34
rect 407 3 410 23
rect 454 3 457 102
rect 516 3 519 39
rect 545 3 548 191
rect 664 180 670 185
rect 582 138 588 143
rect 582 94 585 138
rect 610 73 613 161
rect 617 96 620 141
rect 664 136 667 180
rect 692 115 695 203
rect 699 138 702 183
rect 881 168 884 284
rect 839 165 884 168
rect 774 139 777 150
rect 770 136 783 139
rect 610 3 613 68
rect 692 3 695 110
rect 773 97 776 136
rect 773 94 797 97
rect 802 94 815 97
rect 838 3 841 42
rect 881 3 884 165
rect 7 0 884 3
<< m3contact >>
rect 73 881 78 886
rect 72 770 77 775
rect 84 589 89 594
rect 602 886 607 891
rect 760 727 765 732
rect 76 428 81 433
rect 7 283 12 288
rect 61 255 66 260
rect 771 551 776 556
rect 879 408 884 413
rect 457 283 462 288
rect 265 123 270 128
rect 60 57 65 62
rect 266 3 271 8
rect 771 393 776 398
rect 771 274 776 279
rect 774 150 779 155
<< m123contact >>
rect 317 741 322 746
rect 315 732 320 737
rect 287 652 292 657
rect 279 635 284 640
rect 480 832 485 837
rect 474 740 479 745
rect 583 724 588 729
rect 282 482 287 487
rect 274 462 279 467
rect 300 449 305 454
rect 577 632 582 637
rect 586 611 591 616
rect 431 563 436 568
rect 281 309 286 314
rect 273 296 278 301
rect 388 495 393 500
rect 348 416 353 421
rect 581 552 586 557
rect 496 504 501 509
rect 575 460 580 465
rect 513 408 518 413
rect 283 109 288 114
rect 275 91 280 96
rect 524 216 529 221
rect 586 386 591 391
rect 580 294 585 299
rect 670 215 675 220
rect 588 179 593 184
rect 582 89 587 94
<< metal3 >>
rect 0 920 897 923
rect 0 884 3 920
rect 602 891 605 920
rect 0 881 73 884
rect 0 773 3 881
rect 466 832 480 837
rect 0 770 72 773
rect 0 592 3 770
rect 466 746 470 832
rect 322 741 470 746
rect 474 737 479 740
rect 320 732 479 737
rect 760 732 763 920
rect 569 724 583 728
rect 569 657 573 724
rect 292 653 573 657
rect 284 636 573 639
rect 284 635 577 636
rect 569 632 577 635
rect 531 611 586 614
rect 0 589 84 592
rect 0 431 3 589
rect 436 567 439 568
rect 531 567 534 611
rect 436 564 534 567
rect 436 563 439 564
rect 561 552 581 555
rect 489 504 496 507
rect 489 499 492 504
rect 393 496 492 499
rect 561 487 564 552
rect 894 554 897 920
rect 776 551 897 554
rect 287 484 564 487
rect 279 462 575 465
rect 305 449 325 452
rect 0 428 76 431
rect 0 258 3 428
rect 322 420 325 449
rect 322 417 348 420
rect 875 411 879 413
rect 518 408 879 411
rect 894 396 897 551
rect 776 393 897 396
rect 565 387 586 390
rect 565 314 568 387
rect 286 311 568 314
rect 278 296 580 299
rect 12 283 457 286
rect 894 277 897 393
rect 776 274 897 277
rect 0 255 61 258
rect 0 60 3 255
rect 529 216 670 219
rect 572 179 588 182
rect 0 57 60 60
rect 267 8 270 123
rect 572 114 575 179
rect 894 153 897 274
rect 779 150 897 153
rect 288 111 575 114
rect 280 91 582 94
<< metal4 >>
rect 374 740 377 746
<< labels >>
rlabel metal1 389 711 389 711 7 c1
rlabel metal1 355 710 355 710 3 g0_bar
rlabel metal1 342 622 342 622 3 p1_bar
rlabel metal1 342 596 342 596 3 g1_bar
rlabel metal1 456 604 456 604 7 c2
rlabel metal1 329 524 329 524 3 p2_bar
rlabel metal1 528 434 528 434 7 c3
rlabel metal1 524 217 524 217 1 c4
rlabel metal1 355 217 355 217 1 g3_bar
rlabel metal1 335 145 335 145 1 p4_bar
rlabel metal1 325 26 325 26 1 g4_bar
rlabel metal1 539 65 539 65 7 c5
rlabel metal1 288 634 288 634 1 b1
rlabel metal1 282 634 282 634 3 a1
rlabel metal1 328 742 328 742 1 a0
rlabel metal1 328 735 328 735 1 b0
rlabel metal1 325 408 325 408 1 g2_bar
rlabel metal1 283 458 283 458 1 b2
rlabel metal1 277 458 277 458 3 a2
rlabel metal1 330 336 330 336 1 p3_bar
rlabel metal1 283 291 283 291 1 b3
rlabel metal1 276 291 276 291 3 a3
rlabel metal1 284 89 284 89 1 b4
rlabel metal1 278 89 278 89 3 a4
rlabel metal1 546 749 546 749 1 s0
rlabel metal1 647 641 647 641 7 p1
rlabel metal1 722 647 722 647 7 s1
rlabel metal1 642 469 642 469 1 p2
rlabel metal1 647 303 647 303 1 p3
rlabel metal1 733 304 733 304 7 s3
rlabel metal1 648 98 648 98 1 p4
rlabel metal1 729 140 729 140 1 s4
rlabel metal1 732 469 732 469 7 s2
rlabel metal1 689 827 689 827 1 S0_out
rlabel metal1 169 714 169 714 3 B0_in
rlabel metal1 57 654 57 654 3 B1_in
rlabel metal1 157 575 157 575 1 A1_in
rlabel metal1 48 512 48 512 3 B2_in
rlabel metal1 152 413 152 413 1 A2_in
rlabel metal1 32 359 32 359 3 B3_in
rlabel metal1 145 240 145 240 1 A3_in
rlabel metal1 26 129 26 129 3 B4_in
rlabel metal1 139 42 139 42 1 A4_in
rlabel metal1 844 673 844 673 7 S1_out
rlabel metal1 855 495 855 495 7 S2_out
rlabel metal1 858 337 858 337 7 S3_out
rlabel metal1 856 219 856 219 1 S4_out
rlabel metal1 862 96 862 96 7 COUT_out
rlabel metal1 169 825 169 825 1 A0_in
rlabel metal1 480 899 480 899 5 vdd
rlabel metal2 442 1 442 1 1 gnd
rlabel metal3 480 922 480 922 5 clk
<< end >>
