TSPC D flip flop

.include TSMC_180nm.txt
.param supply=1.8
.param LAMBDA=0.09u
.param width=10*LAMBDA 
.global gnd vdd

Vrail vdd gnd {supply}
Vclk clk gnd pulse 0 1.8 5ns 100ps 100ps 19.9ns 40ns
VD D gnd pulse 0 1.8 0ns 100ps 100ps 34.9ns 70ns

M3 A D vdd vdd CMOSP W={width*4} L={2*LAMBDA}
+ AS={5*4*width*LAMBDA} PS={10*LAMBDA+2*4*width} AD={5*4*width*LAMBDA} PD={10*LAMBDA+2*4*width}

M2 X clk A vdd CMOSP W={width*4} L={2*LAMBDA}
+ AS={5*4*width*LAMBDA} PS={10*LAMBDA+2*4*width} AD={5*4*width*LAMBDA} PD={10*LAMBDA+2*4*width}

M1 X D gnd gnd CMOSN W={width} L={2*LAMBDA}
+ AS={5*width*LAMBDA} PS={10*LAMBDA+2*width} AD={5*width*LAMBDA} PD={10*LAMBDA+2*width}

M6 Y clk vdd vdd CMOSP W={width*2} L={2*LAMBDA}
+ AS={5*2*width*LAMBDA} PS={10*LAMBDA+2*2*width} AD={5*2*width*LAMBDA} PD={10*LAMBDA+2*2*width}

M5 Y X B gnd CMOSN W={width*4} L={2*LAMBDA}
+ AS={5*4*width*LAMBDA} PS={10*LAMBDA+2*4*width} AD={5*4*width*LAMBDA} PD={10*LAMBDA+2*4*width}

M4 B clk gnd gnd CMOSN W={width*4} L={2*LAMBDA}
+ AS={5*4*width*LAMBDA} PS={10*LAMBDA+2*4*width} AD={5*4*width*LAMBDA} PD={10*LAMBDA+2*4*width}

M9 Q_bar Y vdd vdd CMOSP W={width*2} L={2*LAMBDA}
+ AS={5*2*width*LAMBDA} PS={10*LAMBDA+2*2*width} AD={5*2*width*LAMBDA} PD={10*LAMBDA+2*2*width}

M8 Q_bar clk C gnd CMOSN W={width*2} L={2*LAMBDA}
+ AS={5*2*width*LAMBDA} PS={10*LAMBDA+2*2*width} AD={5*2*width*LAMBDA} PD={10*LAMBDA+2*2*width}

M7 C Y gnd gnd CMOSN W={width*2} L={2*LAMBDA}
+ AS={5*2*width*LAMBDA} PS={10*LAMBDA+2*2*width} AD={5*2*width*LAMBDA} PD={10*LAMBDA+2*2*width}

M11 Q Q_bar vdd vdd CMOSP W={width*2} L={2*LAMBDA}
+ AS={5*2*width*LAMBDA} PS={10*LAMBDA+2*2*width} AD={5*2*width*LAMBDA} PD={10*LAMBDA+2*2*width}

M10 Q Q_bar gnd gnd CMOSN W={width} L={2*LAMBDA}
+ AS={5*width*LAMBDA} PS={10*LAMBDA+2*width} AD={5*width*LAMBDA} PD={10*LAMBDA+2*width}

.tran 0.1n 200n

.measure tran tpcq0 TRIG v(clk) val=0.9 RISE=2 TARG v(Q) val=0.9 FALL=1
.measure tran tpcq1 TRIG v(clk) val=0.9 RISE=3 TARG v(Q) val=0.9 RISE=1
.measure tran tcq param = '(tpcq0+tpcq1)/2'
* tcq = 93.22 ps 

.measure tran tsu1 TRIG v(D) val=0.9 FALL=1 TARG v(X) val=0.9 RISE=1
.measure tran tsu0 TRIG v(D) val=0.9 RISE=2 TARG v(X) val=0.9 FALL=2
.measure tran tsu param = '(tsu1+tsu0)/2'
* tsu = 69.69 ps

.measure tran thold TRIG v(clk) val=0.9 RISE=2 TARG v(Y) val=0.9 FALL=1
* thold = 39.03 ps

.control
run
set color0 = white
set color1 = black
set curplottitle = 'NagamallaSaiAbhinav_2024102037'
plot v(Q) v(D)+2 v(clk)+4
.endc