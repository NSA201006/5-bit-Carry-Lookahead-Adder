2 input OR gate

.include TSMC_180nm.txt
.param supply=1.8
.param LAMBDA=0.09u
.param width=10*LAMBDA 
.global gnd vdd

Vrail vdd gnd {supply}
VA A gnd pulse 0 1.8 0ns 100ps 100ps 50ns 100ns
VB B gnd pulse 0 1.8 0ns 100ps 100ps 100ns 200ns

M1 Y_bar A gnd gnd CMOSN W={width} L={2*LAMBDA}
+ AS={5*width*LAMBDA} PS={10*LAMBDA+2*width} AD={5*width*LAMBDA} PD={10*LAMBDA+2*width}

M2 Y_bar B gnd gnd CMOSN W={width} L={2*LAMBDA}
+ AS={5*width*LAMBDA} PS={10*LAMBDA+2*width} AD={5*width*LAMBDA} PD={10*LAMBDA+2*width}

M3 Y_bar A inter vdd CMOSP W={4*width} L={2*LAMBDA}
+ AS={5*4*width*LAMBDA} PS={10*LAMBDA+2*4*width} AD={5*4*width*LAMBDA} PD={10*LAMBDA+2*4*width}

M4 inter B vdd vdd CMOSP W={4*width} L={2*LAMBDA}
+ AS={5*4*width*LAMBDA} PS={10*LAMBDA+2*4*width} AD={5*4*width*LAMBDA} PD={10*LAMBDA+2*4*width}

M5 Y Y_bar vdd vdd CMOSP W={2*width} L={2*LAMBDA}
+ AS={5*2*width*LAMBDA} PS={10*LAMBDA+2*2*width} AD={5*2*width*LAMBDA} PD={10*LAMBDA+2*2*width}

M6 Y Y_bar gnd gnd CMOSN W={width} L={2*LAMBDA}
+ AS={5*width*LAMBDA} PS={10*LAMBDA+2*width} AD={5*width*LAMBDA} PD={10*LAMBDA+2*width}

.tran 0.1n 200n

.control
run
set color0 = white
set color1 = black
set curplottitle = 'NagamallaSaiAbhinav_2024102037'
plot v(Y) v(B)+2 v(A)+4
.endc