magic
tech scmos
timestamp 1763205877
<< nwell >>
rect 0 83 24 115
rect -10 33 26 53
rect -10 1 50 33
rect 57 -24 91 8
rect -10 -97 26 -45
rect 49 -109 107 -77
rect -20 -155 16 -135
rect -20 -187 40 -155
rect 103 -160 139 -140
rect 54 -211 88 -179
rect 103 -192 163 -160
rect -29 -285 7 -233
rect 93 -304 151 -272
rect -22 -346 14 -326
rect -22 -378 38 -346
rect 54 -403 88 -371
rect 98 -377 134 -357
rect 98 -409 158 -377
rect -22 -476 14 -424
rect 56 -488 114 -456
rect -28 -534 8 -514
rect 114 -529 150 -509
rect -28 -535 32 -534
rect -28 -566 66 -535
rect 114 -561 174 -529
rect 32 -567 66 -566
<< ntransistor >>
rect 11 67 13 77
rect 2 -21 4 -11
rect 12 -21 14 -11
rect 37 -17 39 -7
rect 68 -57 70 -37
rect 78 -57 80 -37
rect 2 -119 4 -109
rect 12 -119 14 -109
rect 60 -142 62 -122
rect 70 -142 72 -122
rect 94 -125 96 -115
rect -8 -209 -6 -199
rect 2 -209 4 -199
rect 27 -205 29 -195
rect 115 -214 117 -204
rect 125 -214 127 -204
rect 150 -210 152 -200
rect 65 -244 67 -224
rect 75 -244 77 -224
rect -17 -307 -15 -297
rect -7 -307 -5 -297
rect 104 -337 106 -317
rect 114 -337 116 -317
rect 138 -320 140 -310
rect -10 -400 -8 -390
rect 0 -400 2 -390
rect 25 -396 27 -386
rect 65 -436 67 -416
rect 75 -436 77 -416
rect 110 -431 112 -421
rect 120 -431 122 -421
rect 145 -427 147 -417
rect -10 -498 -8 -488
rect 0 -498 2 -488
rect 67 -521 69 -501
rect 77 -521 79 -501
rect 101 -504 103 -494
rect -16 -588 -14 -578
rect -6 -588 -4 -578
rect 19 -584 21 -574
rect 43 -600 45 -580
rect 53 -600 55 -580
rect 126 -583 128 -573
rect 136 -583 138 -573
rect 161 -579 163 -569
<< ptransistor >>
rect 11 89 13 109
rect 2 7 4 47
rect 12 7 14 47
rect 37 7 39 27
rect 68 -18 70 2
rect 78 -18 80 2
rect 2 -91 4 -51
rect 12 -91 14 -51
rect 60 -103 62 -83
rect 70 -103 72 -83
rect 94 -103 96 -83
rect -8 -181 -6 -141
rect 2 -181 4 -141
rect 27 -181 29 -161
rect 65 -205 67 -185
rect 75 -205 77 -185
rect 115 -186 117 -146
rect 125 -186 127 -146
rect 150 -186 152 -166
rect -17 -279 -15 -239
rect -7 -279 -5 -239
rect 104 -298 106 -278
rect 114 -298 116 -278
rect 138 -298 140 -278
rect -10 -372 -8 -332
rect 0 -372 2 -332
rect 25 -372 27 -352
rect 65 -397 67 -377
rect 75 -397 77 -377
rect 110 -403 112 -363
rect 120 -403 122 -363
rect 145 -403 147 -383
rect -10 -470 -8 -430
rect 0 -470 2 -430
rect 67 -482 69 -462
rect 77 -482 79 -462
rect 101 -482 103 -462
rect -16 -560 -14 -520
rect -6 -560 -4 -520
rect 19 -560 21 -540
rect 43 -561 45 -541
rect 53 -561 55 -541
rect 126 -555 128 -515
rect 136 -555 138 -515
rect 161 -555 163 -535
<< ndiffusion >>
rect 6 71 11 77
rect 10 67 11 71
rect 13 73 14 77
rect 13 67 18 73
rect -3 -17 2 -11
rect 1 -21 2 -17
rect 4 -15 6 -11
rect 10 -15 12 -11
rect 4 -21 12 -15
rect 14 -17 19 -11
rect 32 -13 37 -7
rect 36 -17 37 -13
rect 39 -11 40 -7
rect 39 -17 44 -11
rect 14 -21 15 -17
rect 63 -53 68 -37
rect 67 -57 68 -53
rect 70 -57 78 -37
rect 80 -41 81 -37
rect 80 -57 85 -41
rect -3 -115 2 -109
rect 1 -119 2 -115
rect 4 -113 6 -109
rect 10 -113 12 -109
rect 4 -119 12 -113
rect 14 -115 19 -109
rect 14 -119 15 -115
rect 89 -121 94 -115
rect 55 -138 60 -122
rect 59 -142 60 -138
rect 62 -142 70 -122
rect 72 -126 73 -122
rect 93 -125 94 -121
rect 96 -119 97 -115
rect 96 -125 101 -119
rect 72 -142 77 -126
rect -13 -205 -8 -199
rect -9 -209 -8 -205
rect -6 -203 -4 -199
rect 0 -203 2 -199
rect -6 -209 2 -203
rect 4 -205 9 -199
rect 22 -201 27 -195
rect 26 -205 27 -201
rect 29 -199 30 -195
rect 29 -205 34 -199
rect 4 -209 5 -205
rect 110 -210 115 -204
rect 114 -214 115 -210
rect 117 -208 119 -204
rect 123 -208 125 -204
rect 117 -214 125 -208
rect 127 -210 132 -204
rect 145 -206 150 -200
rect 149 -210 150 -206
rect 152 -204 153 -200
rect 152 -210 157 -204
rect 127 -214 128 -210
rect 60 -240 65 -224
rect 64 -244 65 -240
rect 67 -244 75 -224
rect 77 -228 78 -224
rect 77 -244 82 -228
rect -22 -303 -17 -297
rect -18 -307 -17 -303
rect -15 -301 -13 -297
rect -9 -301 -7 -297
rect -15 -307 -7 -301
rect -5 -303 0 -297
rect -5 -307 -4 -303
rect 133 -316 138 -310
rect 99 -333 104 -317
rect 103 -337 104 -333
rect 106 -337 114 -317
rect 116 -321 117 -317
rect 137 -320 138 -316
rect 140 -314 141 -310
rect 140 -320 145 -314
rect 116 -337 121 -321
rect -15 -396 -10 -390
rect -11 -400 -10 -396
rect -8 -394 -6 -390
rect -2 -394 0 -390
rect -8 -400 0 -394
rect 2 -396 7 -390
rect 20 -392 25 -386
rect 24 -396 25 -392
rect 27 -390 28 -386
rect 27 -396 32 -390
rect 2 -400 3 -396
rect 60 -432 65 -416
rect 64 -436 65 -432
rect 67 -436 75 -416
rect 77 -420 78 -416
rect 77 -436 82 -420
rect 105 -427 110 -421
rect 109 -431 110 -427
rect 112 -425 114 -421
rect 118 -425 120 -421
rect 112 -431 120 -425
rect 122 -427 127 -421
rect 140 -423 145 -417
rect 144 -427 145 -423
rect 147 -421 148 -417
rect 147 -427 152 -421
rect 122 -431 123 -427
rect -15 -494 -10 -488
rect -11 -498 -10 -494
rect -8 -492 -6 -488
rect -2 -492 0 -488
rect -8 -498 0 -492
rect 2 -494 7 -488
rect 2 -498 3 -494
rect 96 -500 101 -494
rect 62 -517 67 -501
rect 66 -521 67 -517
rect 69 -521 77 -501
rect 79 -505 80 -501
rect 100 -504 101 -500
rect 103 -498 104 -494
rect 103 -504 108 -498
rect 79 -521 84 -505
rect -21 -584 -16 -578
rect -17 -588 -16 -584
rect -14 -582 -12 -578
rect -8 -582 -6 -578
rect -14 -588 -6 -582
rect -4 -584 1 -578
rect 14 -580 19 -574
rect 18 -584 19 -580
rect 21 -578 22 -574
rect 21 -584 26 -578
rect 121 -579 126 -573
rect -4 -588 -3 -584
rect 38 -596 43 -580
rect 42 -600 43 -596
rect 45 -600 53 -580
rect 55 -584 56 -580
rect 125 -583 126 -579
rect 128 -577 130 -573
rect 134 -577 136 -573
rect 128 -583 136 -577
rect 138 -579 143 -573
rect 156 -575 161 -569
rect 160 -579 161 -575
rect 163 -573 164 -569
rect 163 -579 168 -573
rect 138 -583 139 -579
rect 55 -600 60 -584
<< pdiffusion >>
rect 10 105 11 109
rect 6 89 11 105
rect 13 93 18 109
rect 13 89 14 93
rect 1 43 2 47
rect -3 7 2 43
rect 4 7 12 47
rect 14 11 19 47
rect 14 7 15 11
rect 36 23 37 27
rect 32 7 37 23
rect 39 11 44 27
rect 39 7 40 11
rect 67 -2 68 2
rect 63 -18 68 -2
rect 70 -14 78 2
rect 70 -18 72 -14
rect 76 -18 78 -14
rect 80 -2 81 2
rect 80 -18 85 -2
rect 1 -55 2 -51
rect -3 -91 2 -55
rect 4 -91 12 -51
rect 14 -87 19 -51
rect 14 -91 15 -87
rect 59 -87 60 -83
rect 55 -103 60 -87
rect 62 -99 70 -83
rect 62 -103 64 -99
rect 68 -103 70 -99
rect 72 -87 73 -83
rect 72 -103 77 -87
rect 93 -87 94 -83
rect 89 -103 94 -87
rect 96 -99 101 -83
rect 96 -103 97 -99
rect -9 -145 -8 -141
rect -13 -181 -8 -145
rect -6 -181 2 -141
rect 4 -177 9 -141
rect 114 -150 115 -146
rect 4 -181 5 -177
rect 26 -165 27 -161
rect 22 -181 27 -165
rect 29 -177 34 -161
rect 29 -181 30 -177
rect 64 -189 65 -185
rect 60 -205 65 -189
rect 67 -201 75 -185
rect 67 -205 69 -201
rect 73 -205 75 -201
rect 77 -189 78 -185
rect 110 -186 115 -150
rect 117 -186 125 -146
rect 127 -182 132 -146
rect 127 -186 128 -182
rect 149 -170 150 -166
rect 145 -186 150 -170
rect 152 -182 157 -166
rect 152 -186 153 -182
rect 77 -205 82 -189
rect -18 -243 -17 -239
rect -22 -279 -17 -243
rect -15 -279 -7 -239
rect -5 -275 0 -239
rect -5 -279 -4 -275
rect 103 -282 104 -278
rect 99 -298 104 -282
rect 106 -294 114 -278
rect 106 -298 108 -294
rect 112 -298 114 -294
rect 116 -282 117 -278
rect 116 -298 121 -282
rect 137 -282 138 -278
rect 133 -298 138 -282
rect 140 -294 145 -278
rect 140 -298 141 -294
rect -11 -336 -10 -332
rect -15 -372 -10 -336
rect -8 -372 0 -332
rect 2 -368 7 -332
rect 2 -372 3 -368
rect 24 -356 25 -352
rect 20 -372 25 -356
rect 27 -368 32 -352
rect 27 -372 28 -368
rect 109 -367 110 -363
rect 64 -381 65 -377
rect 60 -397 65 -381
rect 67 -393 75 -377
rect 67 -397 69 -393
rect 73 -397 75 -393
rect 77 -381 78 -377
rect 77 -397 82 -381
rect 105 -403 110 -367
rect 112 -403 120 -363
rect 122 -399 127 -363
rect 122 -403 123 -399
rect 144 -387 145 -383
rect 140 -403 145 -387
rect 147 -399 152 -383
rect 147 -403 148 -399
rect -11 -434 -10 -430
rect -15 -470 -10 -434
rect -8 -470 0 -430
rect 2 -466 7 -430
rect 2 -470 3 -466
rect 66 -466 67 -462
rect 62 -482 67 -466
rect 69 -478 77 -462
rect 69 -482 71 -478
rect 75 -482 77 -478
rect 79 -466 80 -462
rect 79 -482 84 -466
rect 100 -466 101 -462
rect 96 -482 101 -466
rect 103 -478 108 -462
rect 103 -482 104 -478
rect -17 -524 -16 -520
rect -21 -560 -16 -524
rect -14 -560 -6 -520
rect -4 -556 1 -520
rect 125 -519 126 -515
rect -4 -560 -3 -556
rect 18 -544 19 -540
rect 14 -560 19 -544
rect 21 -556 26 -540
rect 21 -560 22 -556
rect 42 -545 43 -541
rect 38 -561 43 -545
rect 45 -557 53 -541
rect 45 -561 47 -557
rect 51 -561 53 -557
rect 55 -545 56 -541
rect 55 -561 60 -545
rect 121 -555 126 -519
rect 128 -555 136 -515
rect 138 -551 143 -515
rect 138 -555 139 -551
rect 160 -539 161 -535
rect 156 -555 161 -539
rect 163 -551 168 -535
rect 163 -555 164 -551
<< ndcontact >>
rect 6 67 10 71
rect 14 73 18 77
rect -3 -21 1 -17
rect 6 -15 10 -11
rect 32 -17 36 -13
rect 40 -11 44 -7
rect 15 -21 19 -17
rect 63 -57 67 -53
rect 81 -41 85 -37
rect -3 -119 1 -115
rect 6 -113 10 -109
rect 15 -119 19 -115
rect 55 -142 59 -138
rect 73 -126 77 -122
rect 89 -125 93 -121
rect 97 -119 101 -115
rect -13 -209 -9 -205
rect -4 -203 0 -199
rect 22 -205 26 -201
rect 30 -199 34 -195
rect 5 -209 9 -205
rect 110 -214 114 -210
rect 119 -208 123 -204
rect 145 -210 149 -206
rect 153 -204 157 -200
rect 128 -214 132 -210
rect 60 -244 64 -240
rect 78 -228 82 -224
rect -22 -307 -18 -303
rect -13 -301 -9 -297
rect -4 -307 0 -303
rect 99 -337 103 -333
rect 117 -321 121 -317
rect 133 -320 137 -316
rect 141 -314 145 -310
rect -15 -400 -11 -396
rect -6 -394 -2 -390
rect 20 -396 24 -392
rect 28 -390 32 -386
rect 3 -400 7 -396
rect 60 -436 64 -432
rect 78 -420 82 -416
rect 105 -431 109 -427
rect 114 -425 118 -421
rect 140 -427 144 -423
rect 148 -421 152 -417
rect 123 -431 127 -427
rect -15 -498 -11 -494
rect -6 -492 -2 -488
rect 3 -498 7 -494
rect 62 -521 66 -517
rect 80 -505 84 -501
rect 96 -504 100 -500
rect 104 -498 108 -494
rect -21 -588 -17 -584
rect -12 -582 -8 -578
rect 14 -584 18 -580
rect 22 -578 26 -574
rect -3 -588 1 -584
rect 38 -600 42 -596
rect 56 -584 60 -580
rect 121 -583 125 -579
rect 130 -577 134 -573
rect 156 -579 160 -575
rect 164 -573 168 -569
rect 139 -583 143 -579
<< pdcontact >>
rect 6 105 10 109
rect 14 89 18 93
rect -3 43 1 47
rect 15 7 19 11
rect 32 23 36 27
rect 40 7 44 11
rect 63 -2 67 2
rect 72 -18 76 -14
rect 81 -2 85 2
rect -3 -55 1 -51
rect 15 -91 19 -87
rect 55 -87 59 -83
rect 64 -103 68 -99
rect 73 -87 77 -83
rect 89 -87 93 -83
rect 97 -103 101 -99
rect -13 -145 -9 -141
rect 110 -150 114 -146
rect 5 -181 9 -177
rect 22 -165 26 -161
rect 30 -181 34 -177
rect 60 -189 64 -185
rect 69 -205 73 -201
rect 78 -189 82 -185
rect 128 -186 132 -182
rect 145 -170 149 -166
rect 153 -186 157 -182
rect -22 -243 -18 -239
rect -4 -279 0 -275
rect 99 -282 103 -278
rect 108 -298 112 -294
rect 117 -282 121 -278
rect 133 -282 137 -278
rect 141 -298 145 -294
rect -15 -336 -11 -332
rect 3 -372 7 -368
rect 20 -356 24 -352
rect 28 -372 32 -368
rect 105 -367 109 -363
rect 60 -381 64 -377
rect 69 -397 73 -393
rect 78 -381 82 -377
rect 123 -403 127 -399
rect 140 -387 144 -383
rect 148 -403 152 -399
rect -15 -434 -11 -430
rect 3 -470 7 -466
rect 62 -466 66 -462
rect 71 -482 75 -478
rect 80 -466 84 -462
rect 96 -466 100 -462
rect 104 -482 108 -478
rect -21 -524 -17 -520
rect 121 -519 125 -515
rect -3 -560 1 -556
rect 14 -544 18 -540
rect 22 -560 26 -556
rect 38 -545 42 -541
rect 47 -561 51 -557
rect 56 -545 60 -541
rect 139 -555 143 -551
rect 156 -539 160 -535
rect 164 -555 168 -551
<< polysilicon >>
rect 11 109 13 112
rect 11 77 13 89
rect 11 64 13 67
rect 2 47 4 50
rect 12 47 14 50
rect 37 27 39 30
rect 2 -11 4 7
rect 12 -11 14 7
rect 37 -7 39 7
rect 68 2 70 6
rect 78 2 80 6
rect 37 -20 39 -17
rect 2 -24 4 -21
rect 12 -24 14 -21
rect 68 -37 70 -18
rect 78 -37 80 -18
rect 2 -51 4 -48
rect 12 -51 14 -48
rect 68 -60 70 -57
rect 78 -60 80 -57
rect 60 -83 62 -79
rect 70 -83 72 -79
rect 94 -83 96 -80
rect 2 -109 4 -91
rect 12 -109 14 -91
rect 2 -122 4 -119
rect 12 -122 14 -119
rect 60 -122 62 -103
rect 70 -122 72 -103
rect 94 -115 96 -103
rect -8 -141 -6 -138
rect 2 -141 4 -138
rect 94 -128 96 -125
rect 60 -145 62 -142
rect 70 -145 72 -142
rect 115 -146 117 -143
rect 125 -146 127 -143
rect 27 -161 29 -158
rect -8 -199 -6 -181
rect 2 -199 4 -181
rect 27 -195 29 -181
rect 65 -185 67 -181
rect 75 -185 77 -181
rect 150 -166 152 -163
rect 115 -204 117 -186
rect 125 -204 127 -186
rect 150 -200 152 -186
rect 27 -208 29 -205
rect -8 -212 -6 -209
rect 2 -212 4 -209
rect 65 -224 67 -205
rect 75 -224 77 -205
rect 150 -213 152 -210
rect 115 -217 117 -214
rect 125 -217 127 -214
rect -17 -239 -15 -236
rect -7 -239 -5 -236
rect 65 -247 67 -244
rect 75 -247 77 -244
rect 104 -278 106 -274
rect 114 -278 116 -274
rect 138 -278 140 -275
rect -17 -297 -15 -279
rect -7 -297 -5 -279
rect -17 -310 -15 -307
rect -7 -310 -5 -307
rect 104 -317 106 -298
rect 114 -317 116 -298
rect 138 -310 140 -298
rect -10 -332 -8 -329
rect 0 -332 2 -329
rect 138 -323 140 -320
rect 104 -340 106 -337
rect 114 -340 116 -337
rect 25 -352 27 -349
rect 110 -363 112 -360
rect 120 -363 122 -360
rect -10 -390 -8 -372
rect 0 -390 2 -372
rect 25 -386 27 -372
rect 65 -377 67 -373
rect 75 -377 77 -373
rect 25 -399 27 -396
rect -10 -403 -8 -400
rect 0 -403 2 -400
rect 65 -416 67 -397
rect 75 -416 77 -397
rect 145 -383 147 -380
rect -10 -430 -8 -427
rect 0 -430 2 -427
rect 110 -421 112 -403
rect 120 -421 122 -403
rect 145 -417 147 -403
rect 145 -430 147 -427
rect 110 -434 112 -431
rect 120 -434 122 -431
rect 65 -439 67 -436
rect 75 -439 77 -436
rect 67 -462 69 -458
rect 77 -462 79 -458
rect 101 -462 103 -459
rect -10 -488 -8 -470
rect 0 -488 2 -470
rect -10 -501 -8 -498
rect 0 -501 2 -498
rect 67 -501 69 -482
rect 77 -501 79 -482
rect 101 -494 103 -482
rect -16 -520 -14 -517
rect -6 -520 -4 -517
rect 101 -507 103 -504
rect 126 -515 128 -512
rect 136 -515 138 -512
rect 67 -524 69 -521
rect 77 -524 79 -521
rect 19 -540 21 -537
rect 43 -541 45 -537
rect 53 -541 55 -537
rect -16 -578 -14 -560
rect -6 -578 -4 -560
rect 19 -574 21 -560
rect 161 -535 163 -532
rect 43 -580 45 -561
rect 53 -580 55 -561
rect 126 -573 128 -555
rect 136 -573 138 -555
rect 161 -569 163 -555
rect 19 -587 21 -584
rect -16 -591 -14 -588
rect -6 -591 -4 -588
rect 161 -582 163 -579
rect 126 -586 128 -583
rect 136 -586 138 -583
rect 43 -603 45 -600
rect 53 -603 55 -600
<< polycontact >>
rect 7 78 11 82
rect -2 -10 2 -6
rect 8 -4 12 0
rect 33 -6 37 -2
rect 64 -29 68 -25
rect 74 -36 78 -32
rect -2 -108 2 -104
rect 8 -102 12 -98
rect 56 -114 60 -110
rect 66 -121 70 -117
rect 90 -114 94 -110
rect -12 -198 -8 -194
rect -2 -192 2 -188
rect 23 -194 27 -190
rect 111 -203 115 -199
rect 121 -197 125 -193
rect 146 -199 150 -195
rect 61 -216 65 -212
rect 71 -223 75 -219
rect -21 -296 -17 -292
rect -11 -290 -7 -286
rect 100 -309 104 -305
rect 110 -316 114 -312
rect 134 -309 138 -305
rect -14 -389 -10 -385
rect -4 -383 0 -379
rect 21 -385 25 -381
rect 61 -408 65 -404
rect 71 -415 75 -411
rect 106 -420 110 -416
rect 116 -414 120 -410
rect 141 -416 145 -412
rect -14 -487 -10 -483
rect -4 -481 0 -477
rect 63 -493 67 -489
rect 73 -500 77 -496
rect 97 -493 101 -489
rect -20 -577 -16 -573
rect -10 -571 -6 -567
rect 15 -573 19 -569
rect 39 -572 43 -568
rect 49 -579 53 -575
rect 122 -572 126 -568
rect 132 -566 136 -562
rect 157 -568 161 -564
<< metal1 >>
rect 1 116 11 119
rect 6 109 9 116
rect 15 82 18 89
rect -14 78 7 81
rect 15 79 55 82
rect -10 0 -7 78
rect 15 77 18 79
rect 6 63 9 67
rect 6 60 16 63
rect -3 54 30 57
rect -3 47 0 54
rect 27 37 30 54
rect 27 34 35 37
rect 32 27 35 34
rect -10 -3 8 0
rect 16 -2 19 7
rect 41 -2 44 7
rect 63 9 85 12
rect 63 2 66 9
rect 82 2 85 9
rect 16 -5 33 -2
rect -27 -10 -17 -7
rect -12 -10 -2 -7
rect 16 -7 19 -5
rect 41 -5 50 -2
rect 41 -7 44 -5
rect 7 -10 19 -7
rect 7 -11 10 -10
rect -3 -27 0 -21
rect 16 -27 19 -21
rect 32 -27 35 -17
rect -3 -30 35 -27
rect 47 -26 50 -5
rect 47 -29 64 -26
rect 73 -26 76 -18
rect 73 -29 94 -26
rect -35 -36 74 -33
rect 82 -37 85 -29
rect -5 -42 1 -39
rect -3 -51 0 -42
rect 63 -60 66 -57
rect 62 -63 67 -60
rect 55 -76 92 -73
rect 55 -83 58 -76
rect 74 -83 77 -76
rect 89 -83 92 -76
rect -11 -101 8 -98
rect 16 -100 19 -91
rect 16 -103 27 -100
rect -41 -108 -31 -105
rect -26 -108 -2 -105
rect 16 -105 19 -103
rect 7 -108 19 -105
rect -20 -188 -17 -108
rect 7 -109 10 -108
rect -3 -125 0 -119
rect 16 -125 19 -119
rect 24 -118 27 -103
rect 45 -114 56 -111
rect 65 -111 68 -103
rect 98 -110 101 -103
rect 65 -114 90 -111
rect 98 -113 107 -110
rect 24 -121 66 -118
rect 74 -122 77 -114
rect 98 -115 101 -113
rect -3 -128 19 -125
rect -13 -134 20 -131
rect -13 -141 -10 -134
rect 17 -151 20 -134
rect 55 -145 58 -142
rect 89 -145 92 -125
rect 54 -148 92 -145
rect 17 -154 25 -151
rect 22 -161 25 -154
rect -20 -191 -2 -188
rect 6 -190 9 -181
rect 31 -190 34 -181
rect 60 -178 82 -175
rect 60 -185 63 -178
rect 79 -185 82 -178
rect 6 -193 23 -190
rect -33 -198 -12 -195
rect 6 -195 9 -193
rect 31 -193 40 -190
rect 104 -193 107 -113
rect 110 -139 143 -136
rect 110 -146 113 -139
rect 140 -156 143 -139
rect 140 -159 148 -156
rect 145 -166 148 -159
rect 31 -195 34 -193
rect -3 -198 9 -195
rect -3 -199 0 -198
rect -13 -215 -10 -209
rect 6 -215 9 -209
rect 22 -215 25 -205
rect -13 -218 25 -215
rect 37 -213 40 -193
rect 103 -196 121 -193
rect 129 -195 132 -186
rect 154 -195 157 -186
rect 129 -198 146 -195
rect 37 -216 61 -213
rect 70 -213 73 -205
rect 99 -203 111 -200
rect 129 -200 132 -198
rect 154 -198 163 -195
rect 154 -200 157 -198
rect 120 -203 132 -200
rect 99 -213 102 -203
rect 120 -204 123 -203
rect 70 -216 102 -213
rect -29 -224 -22 -221
rect 53 -221 71 -220
rect -17 -223 71 -221
rect -17 -224 56 -223
rect 79 -224 82 -216
rect 110 -220 113 -214
rect 129 -220 132 -214
rect 145 -220 148 -210
rect 110 -223 148 -220
rect -24 -230 -18 -227
rect -22 -239 -19 -230
rect 60 -247 63 -244
rect 59 -250 64 -247
rect 99 -271 136 -268
rect -30 -289 -11 -286
rect -3 -288 0 -279
rect 99 -278 102 -271
rect 118 -278 121 -271
rect 133 -278 136 -271
rect -3 -291 50 -288
rect -55 -296 -21 -293
rect -3 -293 0 -291
rect -12 -296 0 -293
rect -34 -386 -31 -296
rect -12 -297 -9 -296
rect -22 -313 -19 -307
rect -3 -313 0 -307
rect -22 -316 0 -313
rect 47 -313 50 -291
rect 91 -309 100 -306
rect 109 -306 112 -298
rect 142 -305 145 -298
rect 109 -309 134 -306
rect 142 -308 151 -305
rect 47 -316 110 -313
rect 118 -317 121 -309
rect 142 -310 145 -308
rect -15 -325 18 -322
rect -15 -332 -12 -325
rect 15 -342 18 -325
rect 99 -340 102 -337
rect 133 -340 136 -320
rect 15 -345 23 -342
rect 98 -343 136 -340
rect 20 -352 23 -345
rect 148 -346 151 -308
rect 99 -349 151 -346
rect -23 -382 -4 -379
rect 4 -381 7 -372
rect 29 -381 32 -372
rect 60 -370 82 -367
rect 60 -377 63 -370
rect 79 -377 82 -370
rect 4 -384 21 -381
rect -34 -389 -14 -386
rect 4 -386 7 -384
rect 29 -384 38 -381
rect 29 -386 32 -384
rect -5 -389 7 -386
rect -34 -477 -31 -389
rect -5 -390 -2 -389
rect -15 -406 -12 -400
rect 4 -406 7 -400
rect 20 -406 23 -396
rect -15 -409 23 -406
rect 35 -405 38 -384
rect 35 -408 61 -405
rect 70 -405 73 -397
rect 70 -408 88 -405
rect -22 -415 71 -412
rect 79 -416 82 -408
rect -17 -421 -11 -418
rect 85 -417 88 -408
rect 99 -410 102 -349
rect 105 -356 138 -353
rect 105 -363 108 -356
rect 135 -373 138 -356
rect 135 -376 143 -373
rect 140 -383 143 -376
rect 99 -413 116 -410
rect 124 -412 127 -403
rect 149 -412 152 -403
rect 124 -415 141 -412
rect 85 -420 106 -417
rect 124 -417 127 -415
rect 149 -415 158 -412
rect 149 -417 152 -415
rect 115 -420 127 -417
rect 115 -421 118 -420
rect -15 -430 -12 -421
rect 60 -439 63 -436
rect 105 -437 108 -431
rect 124 -437 127 -431
rect 140 -437 143 -427
rect 59 -442 64 -439
rect 105 -440 143 -437
rect 62 -455 99 -452
rect 62 -462 65 -455
rect 81 -462 84 -455
rect 96 -462 99 -455
rect -34 -480 -4 -477
rect 4 -479 7 -470
rect 4 -482 39 -479
rect -34 -487 -14 -484
rect 4 -484 7 -482
rect -5 -487 7 -484
rect -34 -551 -31 -487
rect -5 -488 -2 -487
rect -15 -504 -12 -498
rect 4 -504 7 -498
rect 36 -497 39 -482
rect 55 -493 63 -490
rect 72 -490 75 -482
rect 105 -489 108 -482
rect 72 -493 97 -490
rect 105 -492 114 -489
rect 36 -500 73 -497
rect 81 -501 84 -493
rect 105 -494 108 -492
rect -15 -507 7 -504
rect -21 -513 12 -510
rect -21 -520 -18 -513
rect 9 -530 12 -513
rect 62 -524 65 -521
rect 96 -524 99 -504
rect 61 -527 99 -524
rect 9 -533 17 -530
rect 14 -540 17 -533
rect 38 -534 60 -531
rect 38 -541 41 -534
rect 57 -541 60 -534
rect -42 -554 -31 -551
rect -42 -574 -39 -554
rect -30 -570 -10 -567
rect -2 -569 1 -560
rect 23 -569 26 -560
rect -2 -572 15 -569
rect -42 -577 -20 -574
rect -2 -574 1 -572
rect 23 -572 39 -569
rect 48 -569 51 -561
rect 111 -562 114 -492
rect 121 -508 154 -505
rect 121 -515 124 -508
rect 151 -525 154 -508
rect 151 -528 159 -525
rect 156 -535 159 -528
rect 111 -565 132 -562
rect 140 -564 143 -555
rect 165 -564 168 -555
rect 140 -567 157 -564
rect 48 -572 122 -569
rect 140 -569 143 -567
rect 165 -567 174 -564
rect 165 -569 168 -567
rect 131 -572 143 -569
rect 23 -574 26 -572
rect -11 -577 1 -574
rect -11 -578 -8 -577
rect 29 -579 49 -576
rect -21 -594 -18 -588
rect -2 -594 1 -588
rect 14 -594 17 -584
rect -21 -597 17 -594
rect 29 -603 32 -579
rect 57 -580 60 -572
rect 131 -573 134 -572
rect 121 -589 124 -583
rect 140 -589 143 -583
rect 156 -589 159 -579
rect 121 -592 159 -589
rect 38 -603 41 -600
rect -44 -606 32 -603
rect 37 -606 42 -603
<< m2contact >>
rect 55 79 60 84
rect -17 -12 -12 -7
rect 94 -29 99 -24
rect -40 -38 -35 -33
rect -16 -101 -11 -96
rect -31 -108 -26 -103
rect -38 -198 -33 -193
rect 163 -198 168 -193
rect -22 -224 -17 -219
rect -35 -289 -30 -284
rect 86 -309 91 -304
rect -28 -382 -23 -377
rect -28 -415 -22 -409
rect 50 -493 55 -488
rect -35 -570 -30 -565
<< psm12contact >>
rect 40 -114 45 -109
<< metal2 >>
rect -38 -193 -35 -38
rect -15 -96 -12 -12
rect 55 -99 58 79
rect 40 -102 58 -99
rect -29 -279 -26 -108
rect 40 -109 43 -102
rect -35 -282 -26 -279
rect -35 -284 -29 -282
rect -20 -374 -17 -224
rect 96 -297 99 -29
rect 88 -300 99 -297
rect 88 -304 91 -300
rect -28 -377 -17 -374
rect -28 -555 -25 -415
rect 165 -446 168 -198
rect 50 -449 168 -446
rect 50 -488 53 -449
rect -33 -558 -25 -555
rect -33 -565 -30 -558
<< labels >>
rlabel metal1 5 118 5 118 4 vdd
rlabel metal1 12 61 12 61 1 gnd
rlabel metal1 21 80 21 80 7 c1
rlabel metal1 7 -29 7 -29 1 gnd
rlabel metal1 12 55 12 55 5 vdd
rlabel metal1 -13 79 -13 79 3 g0_bar
rlabel metal1 -26 -9 -26 -9 3 p1_bar
rlabel metal1 74 10 74 10 5 vdd
rlabel metal1 65 -62 65 -62 1 gnd
rlabel metal1 -26 -35 -26 -35 3 g1_bar
rlabel metal1 88 -27 88 -27 7 c2
rlabel metal1 -2 -40 -2 -40 5 vdd
rlabel metal1 7 -127 7 -127 1 gnd
rlabel metal1 -39 -107 -39 -107 3 p2_bar
rlabel metal1 -3 -217 -3 -217 1 gnd
rlabel metal1 2 -133 2 -133 5 vdd
rlabel metal1 70 -74 70 -74 1 vdd
rlabel metal1 75 -147 75 -147 1 gnd
rlabel metal1 62 -249 62 -249 1 gnd
rlabel metal1 71 -177 71 -177 5 vdd
rlabel metal1 -26 -223 -26 -223 1 g2_bar
rlabel metal1 125 -137 125 -137 1 vdd
rlabel metal1 126 -222 126 -222 1 gnd
rlabel metal1 -22 -229 -22 -229 1 vdd
rlabel metal1 -13 -315 -13 -315 1 gnd
rlabel metal1 -51 -295 -51 -295 3 p3_bar
rlabel metal1 -2 -324 -2 -324 1 vdd
rlabel metal1 3 -408 3 -408 1 gnd
rlabel metal1 70 -369 70 -369 1 vdd
rlabel metal1 62 -441 62 -441 1 gnd
rlabel metal1 160 -197 160 -197 7 c3
rlabel metal1 114 -269 114 -269 1 vdd
rlabel metal1 119 -341 119 -341 1 gnd
rlabel metal1 124 -439 124 -439 1 gnd
rlabel metal1 122 -355 122 -355 1 vdd
rlabel metal1 156 -414 156 -414 1 c4
rlabel metal1 -13 -414 -13 -414 1 g3_bar
rlabel metal1 -15 -420 -15 -420 1 vdd
rlabel metal1 -7 -506 -7 -506 1 gnd
rlabel metal1 -33 -486 -33 -486 1 p4_bar
rlabel metal1 -6 -512 -6 -512 1 vdd
rlabel metal1 -1 -596 -1 -596 1 gnd
rlabel metal1 -43 -605 -43 -605 1 g4_bar
rlabel metal1 78 -454 78 -454 1 vdd
rlabel metal1 80 -526 80 -526 1 gnd
rlabel metal1 38 -605 38 -605 1 gnd
rlabel metal1 49 -533 49 -533 1 vdd
rlabel metal1 141 -591 141 -591 1 gnd
rlabel metal1 137 -507 137 -507 1 vdd
rlabel metal1 171 -566 171 -566 7 c5
<< end >>
