magic
tech scmos
timestamp 1763316456
<< nwell >>
rect 214 820 238 852
rect 52 729 86 761
rect 204 730 228 762
rect 244 736 268 768
rect 15 652 49 704
rect 93 697 117 729
rect 317 712 341 744
rect 396 718 420 750
rect 83 647 119 667
rect 83 615 143 647
rect 307 622 331 654
rect 347 628 371 660
rect 386 628 410 660
rect 426 634 450 666
rect 150 590 184 622
rect 15 552 49 584
rect 10 478 44 530
rect 83 517 119 569
rect 315 540 339 572
rect 406 540 430 572
rect 142 505 200 537
rect 73 459 109 479
rect 73 427 133 459
rect 196 454 232 474
rect 10 378 44 410
rect 147 403 181 435
rect 196 422 256 454
rect 305 450 329 482
rect 345 456 369 488
rect 396 450 420 482
rect 436 456 460 488
rect 9 305 43 357
rect 64 329 100 381
rect 320 374 344 406
rect 407 374 431 406
rect 186 310 244 342
rect 71 268 107 288
rect 310 284 334 316
rect 350 290 374 322
rect 397 284 421 316
rect 437 290 461 322
rect 9 205 43 237
rect 71 236 131 268
rect 147 211 181 243
rect 191 237 227 257
rect 191 205 251 237
rect 404 211 428 243
rect 11 105 45 157
rect 71 138 107 190
rect 322 169 346 201
rect 149 126 207 158
rect 394 121 418 153
rect 434 127 458 159
rect 65 80 101 100
rect 207 85 243 105
rect 65 79 125 80
rect 65 48 159 79
rect 207 53 267 85
rect 312 79 336 111
rect 352 85 376 117
rect 125 47 159 48
rect 11 5 45 37
<< ntransistor >>
rect 225 804 227 814
rect 211 772 213 792
rect 240 775 242 795
rect 63 696 65 716
rect 73 696 75 716
rect 215 714 217 724
rect 255 710 257 730
rect 328 696 330 706
rect 407 702 409 712
rect 104 681 106 691
rect 314 664 316 684
rect 343 667 345 687
rect 393 670 395 690
rect 422 673 424 693
rect 26 629 28 639
rect 36 629 38 639
rect 26 598 28 618
rect 36 598 38 618
rect 95 593 97 603
rect 105 593 107 603
rect 130 597 132 607
rect 318 606 320 616
rect 358 602 360 622
rect 397 612 399 622
rect 437 608 439 628
rect 161 557 163 577
rect 171 557 173 577
rect 326 524 328 534
rect 417 524 419 534
rect 95 495 97 505
rect 105 495 107 505
rect 21 455 23 465
rect 31 455 33 465
rect 21 424 23 444
rect 31 424 33 444
rect 153 472 155 492
rect 163 472 165 492
rect 187 489 189 499
rect 312 492 314 512
rect 341 495 343 515
rect 403 492 405 512
rect 432 495 434 515
rect 85 405 87 415
rect 95 405 97 415
rect 120 409 122 419
rect 316 434 318 444
rect 356 430 358 450
rect 407 434 409 444
rect 447 430 449 450
rect 208 400 210 410
rect 218 400 220 410
rect 243 404 245 414
rect 158 370 160 390
rect 168 370 170 390
rect 331 358 333 368
rect 418 358 420 368
rect 76 307 78 317
rect 86 307 88 317
rect 317 326 319 346
rect 346 329 348 349
rect 404 326 406 346
rect 433 329 435 349
rect 20 282 22 292
rect 30 282 32 292
rect 20 251 22 271
rect 30 251 32 271
rect 197 277 199 297
rect 207 277 209 297
rect 231 294 233 304
rect 321 268 323 278
rect 361 264 363 284
rect 408 268 410 278
rect 448 264 450 284
rect 83 214 85 224
rect 93 214 95 224
rect 118 218 120 228
rect 158 178 160 198
rect 168 178 170 198
rect 203 183 205 193
rect 213 183 215 193
rect 238 187 240 197
rect 415 195 417 205
rect 401 163 403 183
rect 430 166 432 186
rect 333 153 335 163
rect 83 116 85 126
rect 93 116 95 126
rect 319 121 321 141
rect 348 124 350 144
rect 22 82 24 92
rect 32 82 34 92
rect 22 51 24 71
rect 32 51 34 71
rect 160 93 162 113
rect 170 93 172 113
rect 194 110 196 120
rect 405 105 407 115
rect 445 101 447 121
rect 323 63 325 73
rect 363 59 365 79
rect 77 26 79 36
rect 87 26 89 36
rect 112 30 114 40
rect 136 14 138 34
rect 146 14 148 34
rect 219 31 221 41
rect 229 31 231 41
rect 254 35 256 45
<< ptransistor >>
rect 225 826 227 846
rect 63 735 65 755
rect 73 735 75 755
rect 215 736 217 756
rect 255 742 257 762
rect 26 658 28 698
rect 36 658 38 698
rect 104 703 106 723
rect 328 718 330 738
rect 407 724 409 744
rect 95 621 97 661
rect 105 621 107 661
rect 130 621 132 641
rect 318 628 320 648
rect 358 634 360 654
rect 397 634 399 654
rect 437 640 439 660
rect 161 596 163 616
rect 171 596 173 616
rect 26 558 28 578
rect 36 558 38 578
rect 21 484 23 524
rect 31 484 33 524
rect 95 523 97 563
rect 105 523 107 563
rect 326 546 328 566
rect 417 546 419 566
rect 153 511 155 531
rect 163 511 165 531
rect 187 511 189 531
rect 85 433 87 473
rect 95 433 97 473
rect 120 433 122 453
rect 158 409 160 429
rect 168 409 170 429
rect 208 428 210 468
rect 218 428 220 468
rect 316 456 318 476
rect 356 462 358 482
rect 243 428 245 448
rect 407 456 409 476
rect 447 462 449 482
rect 21 384 23 404
rect 31 384 33 404
rect 20 311 22 351
rect 30 311 32 351
rect 76 335 78 375
rect 86 335 88 375
rect 331 380 333 400
rect 418 380 420 400
rect 197 316 199 336
rect 207 316 209 336
rect 231 316 233 336
rect 83 242 85 282
rect 93 242 95 282
rect 321 290 323 310
rect 361 296 363 316
rect 408 290 410 310
rect 448 296 450 316
rect 118 242 120 262
rect 20 211 22 231
rect 30 211 32 231
rect 158 217 160 237
rect 168 217 170 237
rect 203 211 205 251
rect 213 211 215 251
rect 238 211 240 231
rect 415 217 417 237
rect 22 111 24 151
rect 32 111 34 151
rect 83 144 85 184
rect 93 144 95 184
rect 333 175 335 195
rect 160 132 162 152
rect 170 132 172 152
rect 194 132 196 152
rect 405 127 407 147
rect 445 133 447 153
rect 77 54 79 94
rect 87 54 89 94
rect 112 54 114 74
rect 136 53 138 73
rect 146 53 148 73
rect 219 59 221 99
rect 229 59 231 99
rect 323 85 325 105
rect 363 91 365 111
rect 254 59 256 79
rect 22 11 24 31
rect 32 11 34 31
<< ndiffusion >>
rect 220 808 225 814
rect 224 804 225 808
rect 227 810 228 814
rect 227 804 232 810
rect 205 777 211 792
rect 210 772 211 777
rect 213 776 218 792
rect 213 772 214 776
rect 234 780 240 795
rect 239 775 240 780
rect 242 779 247 795
rect 242 775 243 779
rect 58 700 63 716
rect 62 696 63 700
rect 65 696 73 716
rect 75 712 76 716
rect 75 696 80 712
rect 210 718 215 724
rect 214 714 215 718
rect 217 720 218 724
rect 217 714 222 720
rect 250 714 255 730
rect 254 710 255 714
rect 257 726 258 730
rect 257 710 262 726
rect 402 706 407 712
rect 323 700 328 706
rect 327 696 328 700
rect 330 702 331 706
rect 406 702 407 706
rect 409 708 410 712
rect 409 702 414 708
rect 330 696 335 702
rect 99 685 104 691
rect 103 681 104 685
rect 106 687 107 691
rect 106 681 111 687
rect 308 669 314 684
rect 313 664 314 669
rect 316 668 321 684
rect 316 664 317 668
rect 337 672 343 687
rect 342 667 343 672
rect 345 671 350 687
rect 345 667 346 671
rect 387 675 393 690
rect 392 670 393 675
rect 395 674 400 690
rect 395 670 396 674
rect 416 678 422 693
rect 421 673 422 678
rect 424 677 429 693
rect 424 673 425 677
rect 21 633 26 639
rect 25 629 26 633
rect 28 635 30 639
rect 34 635 36 639
rect 28 629 36 635
rect 38 633 43 639
rect 38 629 39 633
rect 25 614 26 618
rect 21 598 26 614
rect 28 598 36 618
rect 38 602 43 618
rect 38 598 39 602
rect 90 597 95 603
rect 94 593 95 597
rect 97 599 99 603
rect 103 599 105 603
rect 97 593 105 599
rect 107 597 112 603
rect 125 601 130 607
rect 129 597 130 601
rect 132 603 133 607
rect 132 597 137 603
rect 107 593 108 597
rect 313 610 318 616
rect 317 606 318 610
rect 320 612 321 616
rect 320 606 325 612
rect 353 606 358 622
rect 357 602 358 606
rect 360 618 361 622
rect 360 602 365 618
rect 392 616 397 622
rect 396 612 397 616
rect 399 618 400 622
rect 399 612 404 618
rect 432 612 437 628
rect 436 608 437 612
rect 439 624 440 628
rect 439 608 444 624
rect 156 561 161 577
rect 160 557 161 561
rect 163 557 171 577
rect 173 573 174 577
rect 173 557 178 573
rect 321 528 326 534
rect 325 524 326 528
rect 328 530 329 534
rect 328 524 333 530
rect 412 528 417 534
rect 416 524 417 528
rect 419 530 420 534
rect 419 524 424 530
rect 90 499 95 505
rect 94 495 95 499
rect 97 501 99 505
rect 103 501 105 505
rect 97 495 105 501
rect 107 499 112 505
rect 107 495 108 499
rect 182 493 187 499
rect 148 476 153 492
rect 16 459 21 465
rect 20 455 21 459
rect 23 461 25 465
rect 29 461 31 465
rect 23 455 31 461
rect 33 459 38 465
rect 33 455 34 459
rect 20 440 21 444
rect 16 424 21 440
rect 23 424 31 444
rect 33 428 38 444
rect 152 472 153 476
rect 155 472 163 492
rect 165 488 166 492
rect 186 489 187 493
rect 189 495 190 499
rect 189 489 194 495
rect 306 497 312 512
rect 311 492 312 497
rect 314 496 319 512
rect 314 492 315 496
rect 335 500 341 515
rect 340 495 341 500
rect 343 499 348 515
rect 343 495 344 499
rect 397 497 403 512
rect 402 492 403 497
rect 405 496 410 512
rect 405 492 406 496
rect 426 500 432 515
rect 431 495 432 500
rect 434 499 439 515
rect 434 495 435 499
rect 165 472 170 488
rect 33 424 34 428
rect 80 409 85 415
rect 84 405 85 409
rect 87 411 89 415
rect 93 411 95 415
rect 87 405 95 411
rect 97 409 102 415
rect 115 413 120 419
rect 119 409 120 413
rect 122 415 123 419
rect 122 409 127 415
rect 311 438 316 444
rect 315 434 316 438
rect 318 440 319 444
rect 318 434 323 440
rect 351 434 356 450
rect 355 430 356 434
rect 358 446 359 450
rect 358 430 363 446
rect 402 438 407 444
rect 406 434 407 438
rect 409 440 410 444
rect 409 434 414 440
rect 442 434 447 450
rect 446 430 447 434
rect 449 446 450 450
rect 449 430 454 446
rect 97 405 98 409
rect 203 404 208 410
rect 207 400 208 404
rect 210 406 212 410
rect 216 406 218 410
rect 210 400 218 406
rect 220 404 225 410
rect 238 408 243 414
rect 242 404 243 408
rect 245 410 246 414
rect 245 404 250 410
rect 220 400 221 404
rect 153 374 158 390
rect 157 370 158 374
rect 160 370 168 390
rect 170 386 171 390
rect 170 370 175 386
rect 326 362 331 368
rect 330 358 331 362
rect 333 364 334 368
rect 333 358 338 364
rect 413 362 418 368
rect 417 358 418 362
rect 420 364 421 368
rect 420 358 425 364
rect 71 311 76 317
rect 75 307 76 311
rect 78 313 80 317
rect 84 313 86 317
rect 78 307 86 313
rect 88 311 93 317
rect 311 331 317 346
rect 316 326 317 331
rect 319 330 324 346
rect 319 326 320 330
rect 340 334 346 349
rect 345 329 346 334
rect 348 333 353 349
rect 348 329 349 333
rect 398 331 404 346
rect 403 326 404 331
rect 406 330 411 346
rect 406 326 407 330
rect 427 334 433 349
rect 432 329 433 334
rect 435 333 440 349
rect 435 329 436 333
rect 88 307 89 311
rect 226 298 231 304
rect 15 286 20 292
rect 19 282 20 286
rect 22 288 24 292
rect 28 288 30 292
rect 22 282 30 288
rect 32 286 37 292
rect 32 282 33 286
rect 19 267 20 271
rect 15 251 20 267
rect 22 251 30 271
rect 32 255 37 271
rect 32 251 33 255
rect 192 281 197 297
rect 196 277 197 281
rect 199 277 207 297
rect 209 293 210 297
rect 230 294 231 298
rect 233 300 234 304
rect 233 294 238 300
rect 209 277 214 293
rect 316 272 321 278
rect 320 268 321 272
rect 323 274 324 278
rect 323 268 328 274
rect 356 268 361 284
rect 360 264 361 268
rect 363 280 364 284
rect 363 264 368 280
rect 403 272 408 278
rect 407 268 408 272
rect 410 274 411 278
rect 410 268 415 274
rect 443 268 448 284
rect 447 264 448 268
rect 450 280 451 284
rect 450 264 455 280
rect 78 218 83 224
rect 82 214 83 218
rect 85 220 87 224
rect 91 220 93 224
rect 85 214 93 220
rect 95 218 100 224
rect 113 222 118 228
rect 117 218 118 222
rect 120 224 121 228
rect 120 218 125 224
rect 95 214 96 218
rect 153 182 158 198
rect 157 178 158 182
rect 160 178 168 198
rect 170 194 171 198
rect 170 178 175 194
rect 410 199 415 205
rect 198 187 203 193
rect 202 183 203 187
rect 205 189 207 193
rect 211 189 213 193
rect 205 183 213 189
rect 215 187 220 193
rect 233 191 238 197
rect 237 187 238 191
rect 240 193 241 197
rect 414 195 415 199
rect 417 201 418 205
rect 417 195 422 201
rect 240 187 245 193
rect 215 183 216 187
rect 395 168 401 183
rect 400 163 401 168
rect 403 167 408 183
rect 403 163 404 167
rect 424 171 430 186
rect 429 166 430 171
rect 432 170 437 186
rect 432 166 433 170
rect 328 157 333 163
rect 332 153 333 157
rect 335 159 336 163
rect 335 153 340 159
rect 78 120 83 126
rect 82 116 83 120
rect 85 122 87 126
rect 91 122 93 126
rect 85 116 93 122
rect 95 120 100 126
rect 95 116 96 120
rect 313 126 319 141
rect 318 121 319 126
rect 321 125 326 141
rect 321 121 322 125
rect 342 129 348 144
rect 347 124 348 129
rect 350 128 355 144
rect 350 124 351 128
rect 189 114 194 120
rect 155 97 160 113
rect 17 86 22 92
rect 21 82 22 86
rect 24 88 26 92
rect 30 88 32 92
rect 24 82 32 88
rect 34 86 39 92
rect 34 82 35 86
rect 21 67 22 71
rect 17 51 22 67
rect 24 51 32 71
rect 34 55 39 71
rect 34 51 35 55
rect 159 93 160 97
rect 162 93 170 113
rect 172 109 173 113
rect 193 110 194 114
rect 196 116 197 120
rect 196 110 201 116
rect 172 93 177 109
rect 400 109 405 115
rect 404 105 405 109
rect 407 111 408 115
rect 407 105 412 111
rect 440 105 445 121
rect 444 101 445 105
rect 447 117 448 121
rect 447 101 452 117
rect 318 67 323 73
rect 322 63 323 67
rect 325 69 326 73
rect 325 63 330 69
rect 358 63 363 79
rect 362 59 363 63
rect 365 75 366 79
rect 365 59 370 75
rect 72 30 77 36
rect 76 26 77 30
rect 79 32 81 36
rect 85 32 87 36
rect 79 26 87 32
rect 89 30 94 36
rect 107 34 112 40
rect 111 30 112 34
rect 114 36 115 40
rect 114 30 119 36
rect 214 35 219 41
rect 89 26 90 30
rect 131 18 136 34
rect 135 14 136 18
rect 138 14 146 34
rect 148 30 149 34
rect 218 31 219 35
rect 221 37 223 41
rect 227 37 229 41
rect 221 31 229 37
rect 231 35 236 41
rect 249 39 254 45
rect 253 35 254 39
rect 256 41 257 45
rect 256 35 261 41
rect 231 31 232 35
rect 148 14 153 30
<< pdiffusion >>
rect 224 842 225 846
rect 220 826 225 842
rect 227 830 232 846
rect 227 826 228 830
rect 254 758 255 762
rect 62 751 63 755
rect 58 735 63 751
rect 65 739 73 755
rect 65 735 67 739
rect 71 735 73 739
rect 75 751 76 755
rect 75 735 80 751
rect 214 752 215 756
rect 210 736 215 752
rect 217 740 222 756
rect 250 742 255 758
rect 257 746 262 762
rect 257 742 258 746
rect 217 736 218 740
rect 406 740 407 744
rect 327 734 328 738
rect 103 719 104 723
rect 25 694 26 698
rect 21 658 26 694
rect 28 658 36 698
rect 38 662 43 698
rect 99 703 104 719
rect 106 707 111 723
rect 323 718 328 734
rect 330 722 335 738
rect 402 724 407 740
rect 409 728 414 744
rect 409 724 410 728
rect 330 718 331 722
rect 106 703 107 707
rect 38 658 39 662
rect 94 657 95 661
rect 90 621 95 657
rect 97 621 105 661
rect 107 625 112 661
rect 436 656 437 660
rect 357 650 358 654
rect 317 644 318 648
rect 107 621 108 625
rect 129 637 130 641
rect 125 621 130 637
rect 132 625 137 641
rect 313 628 318 644
rect 320 632 325 648
rect 353 634 358 650
rect 360 638 365 654
rect 360 634 361 638
rect 396 650 397 654
rect 392 634 397 650
rect 399 638 404 654
rect 432 640 437 656
rect 439 644 444 660
rect 439 640 440 644
rect 399 634 400 638
rect 320 628 321 632
rect 132 621 133 625
rect 160 612 161 616
rect 156 596 161 612
rect 163 600 171 616
rect 163 596 165 600
rect 169 596 171 600
rect 173 612 174 616
rect 173 596 178 612
rect 21 562 26 578
rect 25 558 26 562
rect 28 574 30 578
rect 34 574 36 578
rect 28 558 36 574
rect 38 562 43 578
rect 38 558 39 562
rect 94 559 95 563
rect 20 520 21 524
rect 16 484 21 520
rect 23 484 31 524
rect 33 488 38 524
rect 90 523 95 559
rect 97 523 105 563
rect 107 527 112 563
rect 325 562 326 566
rect 321 546 326 562
rect 328 550 333 566
rect 328 546 329 550
rect 416 562 417 566
rect 412 546 417 562
rect 419 550 424 566
rect 419 546 420 550
rect 107 523 108 527
rect 152 527 153 531
rect 148 511 153 527
rect 155 515 163 531
rect 155 511 157 515
rect 161 511 163 515
rect 165 527 166 531
rect 165 511 170 527
rect 186 527 187 531
rect 182 511 187 527
rect 189 515 194 531
rect 189 511 190 515
rect 33 484 34 488
rect 84 469 85 473
rect 80 433 85 469
rect 87 433 95 473
rect 97 437 102 473
rect 355 478 356 482
rect 315 472 316 476
rect 207 464 208 468
rect 97 433 98 437
rect 119 449 120 453
rect 115 433 120 449
rect 122 437 127 453
rect 122 433 123 437
rect 157 425 158 429
rect 153 409 158 425
rect 160 413 168 429
rect 160 409 162 413
rect 166 409 168 413
rect 170 425 171 429
rect 203 428 208 464
rect 210 428 218 468
rect 220 432 225 468
rect 311 456 316 472
rect 318 460 323 476
rect 351 462 356 478
rect 358 466 363 482
rect 446 478 447 482
rect 358 462 359 466
rect 406 472 407 476
rect 318 456 319 460
rect 220 428 221 432
rect 242 444 243 448
rect 238 428 243 444
rect 245 432 250 448
rect 402 456 407 472
rect 409 460 414 476
rect 442 462 447 478
rect 449 466 454 482
rect 449 462 450 466
rect 409 456 410 460
rect 245 428 246 432
rect 170 409 175 425
rect 16 388 21 404
rect 20 384 21 388
rect 23 400 25 404
rect 29 400 31 404
rect 23 384 31 400
rect 33 388 38 404
rect 330 396 331 400
rect 33 384 34 388
rect 75 371 76 375
rect 19 347 20 351
rect 15 311 20 347
rect 22 311 30 351
rect 32 315 37 351
rect 71 335 76 371
rect 78 335 86 375
rect 88 339 93 375
rect 326 380 331 396
rect 333 384 338 400
rect 333 380 334 384
rect 417 396 418 400
rect 413 380 418 396
rect 420 384 425 400
rect 420 380 421 384
rect 88 335 89 339
rect 196 332 197 336
rect 32 311 33 315
rect 192 316 197 332
rect 199 320 207 336
rect 199 316 201 320
rect 205 316 207 320
rect 209 332 210 336
rect 209 316 214 332
rect 230 332 231 336
rect 226 316 231 332
rect 233 320 238 336
rect 233 316 234 320
rect 360 312 361 316
rect 320 306 321 310
rect 82 278 83 282
rect 78 242 83 278
rect 85 242 93 282
rect 95 246 100 282
rect 316 290 321 306
rect 323 294 328 310
rect 356 296 361 312
rect 363 300 368 316
rect 447 312 448 316
rect 363 296 364 300
rect 407 306 408 310
rect 323 290 324 294
rect 403 290 408 306
rect 410 294 415 310
rect 443 296 448 312
rect 450 300 455 316
rect 450 296 451 300
rect 410 290 411 294
rect 95 242 96 246
rect 117 258 118 262
rect 113 242 118 258
rect 120 246 125 262
rect 120 242 121 246
rect 202 247 203 251
rect 15 215 20 231
rect 19 211 20 215
rect 22 227 24 231
rect 28 227 30 231
rect 22 211 30 227
rect 32 215 37 231
rect 157 233 158 237
rect 32 211 33 215
rect 153 217 158 233
rect 160 221 168 237
rect 160 217 162 221
rect 166 217 168 221
rect 170 233 171 237
rect 170 217 175 233
rect 198 211 203 247
rect 205 211 213 251
rect 215 215 220 251
rect 414 233 415 237
rect 215 211 216 215
rect 237 227 238 231
rect 233 211 238 227
rect 240 215 245 231
rect 410 217 415 233
rect 417 221 422 237
rect 417 217 418 221
rect 240 211 241 215
rect 82 180 83 184
rect 21 147 22 151
rect 17 111 22 147
rect 24 111 32 151
rect 34 115 39 151
rect 78 144 83 180
rect 85 144 93 184
rect 95 148 100 184
rect 332 191 333 195
rect 328 175 333 191
rect 335 179 340 195
rect 335 175 336 179
rect 95 144 96 148
rect 159 148 160 152
rect 155 132 160 148
rect 162 136 170 152
rect 162 132 164 136
rect 168 132 170 136
rect 172 148 173 152
rect 172 132 177 148
rect 193 148 194 152
rect 189 132 194 148
rect 196 136 201 152
rect 444 149 445 153
rect 196 132 197 136
rect 34 111 35 115
rect 404 143 405 147
rect 400 127 405 143
rect 407 131 412 147
rect 440 133 445 149
rect 447 137 452 153
rect 447 133 448 137
rect 407 127 408 131
rect 76 90 77 94
rect 72 54 77 90
rect 79 54 87 94
rect 89 58 94 94
rect 362 107 363 111
rect 322 101 323 105
rect 218 95 219 99
rect 89 54 90 58
rect 111 70 112 74
rect 107 54 112 70
rect 114 58 119 74
rect 114 54 115 58
rect 135 69 136 73
rect 131 53 136 69
rect 138 57 146 73
rect 138 53 140 57
rect 144 53 146 57
rect 148 69 149 73
rect 148 53 153 69
rect 214 59 219 95
rect 221 59 229 99
rect 231 63 236 99
rect 318 85 323 101
rect 325 89 330 105
rect 358 91 363 107
rect 365 95 370 111
rect 365 91 366 95
rect 325 85 326 89
rect 231 59 232 63
rect 253 75 254 79
rect 249 59 254 75
rect 256 63 261 79
rect 256 59 257 63
rect 17 15 22 31
rect 21 11 22 15
rect 24 27 26 31
rect 30 27 32 31
rect 24 11 32 27
rect 34 15 39 31
rect 34 11 35 15
<< ndcontact >>
rect 220 804 224 808
rect 228 810 232 814
rect 214 772 218 776
rect 243 775 247 779
rect 58 696 62 700
rect 76 712 80 716
rect 210 714 214 718
rect 218 720 222 724
rect 250 710 254 714
rect 258 726 262 730
rect 323 696 327 700
rect 331 702 335 706
rect 402 702 406 706
rect 410 708 414 712
rect 99 681 103 685
rect 107 687 111 691
rect 317 664 321 668
rect 346 667 350 671
rect 396 670 400 674
rect 425 673 429 677
rect 21 629 25 633
rect 30 635 34 639
rect 39 629 43 633
rect 21 614 25 618
rect 39 598 43 602
rect 90 593 94 597
rect 99 599 103 603
rect 125 597 129 601
rect 133 603 137 607
rect 108 593 112 597
rect 313 606 317 610
rect 321 612 325 616
rect 353 602 357 606
rect 361 618 365 622
rect 392 612 396 616
rect 400 618 404 622
rect 432 608 436 612
rect 440 624 444 628
rect 156 557 160 561
rect 174 573 178 577
rect 321 524 325 528
rect 329 530 333 534
rect 412 524 416 528
rect 420 530 424 534
rect 90 495 94 499
rect 99 501 103 505
rect 108 495 112 499
rect 16 455 20 459
rect 25 461 29 465
rect 34 455 38 459
rect 16 440 20 444
rect 148 472 152 476
rect 166 488 170 492
rect 182 489 186 493
rect 190 495 194 499
rect 315 492 319 496
rect 344 495 348 499
rect 406 492 410 496
rect 435 495 439 499
rect 34 424 38 428
rect 80 405 84 409
rect 89 411 93 415
rect 115 409 119 413
rect 123 415 127 419
rect 311 434 315 438
rect 319 440 323 444
rect 351 430 355 434
rect 359 446 363 450
rect 402 434 406 438
rect 410 440 414 444
rect 442 430 446 434
rect 450 446 454 450
rect 98 405 102 409
rect 203 400 207 404
rect 212 406 216 410
rect 238 404 242 408
rect 246 410 250 414
rect 221 400 225 404
rect 153 370 157 374
rect 171 386 175 390
rect 326 358 330 362
rect 334 364 338 368
rect 413 358 417 362
rect 421 364 425 368
rect 71 307 75 311
rect 80 313 84 317
rect 320 326 324 330
rect 349 329 353 333
rect 407 326 411 330
rect 436 329 440 333
rect 89 307 93 311
rect 15 282 19 286
rect 24 288 28 292
rect 33 282 37 286
rect 15 267 19 271
rect 33 251 37 255
rect 192 277 196 281
rect 210 293 214 297
rect 226 294 230 298
rect 234 300 238 304
rect 316 268 320 272
rect 324 274 328 278
rect 356 264 360 268
rect 364 280 368 284
rect 403 268 407 272
rect 411 274 415 278
rect 443 264 447 268
rect 451 280 455 284
rect 78 214 82 218
rect 87 220 91 224
rect 113 218 117 222
rect 121 224 125 228
rect 96 214 100 218
rect 153 178 157 182
rect 171 194 175 198
rect 198 183 202 187
rect 207 189 211 193
rect 233 187 237 191
rect 241 193 245 197
rect 410 195 414 199
rect 418 201 422 205
rect 216 183 220 187
rect 404 163 408 167
rect 433 166 437 170
rect 328 153 332 157
rect 336 159 340 163
rect 78 116 82 120
rect 87 122 91 126
rect 96 116 100 120
rect 322 121 326 125
rect 351 124 355 128
rect 17 82 21 86
rect 26 88 30 92
rect 35 82 39 86
rect 17 67 21 71
rect 35 51 39 55
rect 155 93 159 97
rect 173 109 177 113
rect 189 110 193 114
rect 197 116 201 120
rect 400 105 404 109
rect 408 111 412 115
rect 440 101 444 105
rect 448 117 452 121
rect 318 63 322 67
rect 326 69 330 73
rect 358 59 362 63
rect 366 75 370 79
rect 72 26 76 30
rect 81 32 85 36
rect 107 30 111 34
rect 115 36 119 40
rect 90 26 94 30
rect 131 14 135 18
rect 149 30 153 34
rect 214 31 218 35
rect 223 37 227 41
rect 249 35 253 39
rect 257 41 261 45
rect 232 31 236 35
<< pdcontact >>
rect 220 842 224 846
rect 228 826 232 830
rect 250 758 254 762
rect 58 751 62 755
rect 67 735 71 739
rect 76 751 80 755
rect 210 752 214 756
rect 258 742 262 746
rect 218 736 222 740
rect 402 740 406 744
rect 323 734 327 738
rect 99 719 103 723
rect 21 694 25 698
rect 410 724 414 728
rect 331 718 335 722
rect 107 703 111 707
rect 39 658 43 662
rect 90 657 94 661
rect 432 656 436 660
rect 353 650 357 654
rect 313 644 317 648
rect 108 621 112 625
rect 125 637 129 641
rect 361 634 365 638
rect 392 650 396 654
rect 440 640 444 644
rect 400 634 404 638
rect 321 628 325 632
rect 133 621 137 625
rect 156 612 160 616
rect 165 596 169 600
rect 174 612 178 616
rect 21 558 25 562
rect 30 574 34 578
rect 39 558 43 562
rect 90 559 94 563
rect 16 520 20 524
rect 321 562 325 566
rect 329 546 333 550
rect 412 562 416 566
rect 420 546 424 550
rect 108 523 112 527
rect 148 527 152 531
rect 157 511 161 515
rect 166 527 170 531
rect 182 527 186 531
rect 190 511 194 515
rect 34 484 38 488
rect 80 469 84 473
rect 351 478 355 482
rect 311 472 315 476
rect 203 464 207 468
rect 98 433 102 437
rect 115 449 119 453
rect 123 433 127 437
rect 153 425 157 429
rect 162 409 166 413
rect 171 425 175 429
rect 442 478 446 482
rect 359 462 363 466
rect 402 472 406 476
rect 319 456 323 460
rect 221 428 225 432
rect 238 444 242 448
rect 450 462 454 466
rect 410 456 414 460
rect 246 428 250 432
rect 16 384 20 388
rect 25 400 29 404
rect 326 396 330 400
rect 34 384 38 388
rect 71 371 75 375
rect 15 347 19 351
rect 334 380 338 384
rect 413 396 417 400
rect 421 380 425 384
rect 89 335 93 339
rect 192 332 196 336
rect 33 311 37 315
rect 201 316 205 320
rect 210 332 214 336
rect 226 332 230 336
rect 234 316 238 320
rect 356 312 360 316
rect 316 306 320 310
rect 78 278 82 282
rect 443 312 447 316
rect 364 296 368 300
rect 403 306 407 310
rect 324 290 328 294
rect 451 296 455 300
rect 411 290 415 294
rect 96 242 100 246
rect 113 258 117 262
rect 121 242 125 246
rect 198 247 202 251
rect 15 211 19 215
rect 24 227 28 231
rect 153 233 157 237
rect 33 211 37 215
rect 162 217 166 221
rect 171 233 175 237
rect 410 233 414 237
rect 216 211 220 215
rect 233 227 237 231
rect 418 217 422 221
rect 241 211 245 215
rect 78 180 82 184
rect 17 147 21 151
rect 328 191 332 195
rect 336 175 340 179
rect 96 144 100 148
rect 155 148 159 152
rect 164 132 168 136
rect 173 148 177 152
rect 189 148 193 152
rect 440 149 444 153
rect 197 132 201 136
rect 35 111 39 115
rect 400 143 404 147
rect 448 133 452 137
rect 408 127 412 131
rect 72 90 76 94
rect 358 107 362 111
rect 318 101 322 105
rect 214 95 218 99
rect 90 54 94 58
rect 107 70 111 74
rect 115 54 119 58
rect 131 69 135 73
rect 140 53 144 57
rect 149 69 153 73
rect 366 91 370 95
rect 326 85 330 89
rect 232 59 236 63
rect 249 75 253 79
rect 257 59 261 63
rect 17 11 21 15
rect 26 27 30 31
rect 35 11 39 15
<< polysilicon >>
rect 225 846 227 849
rect 225 814 227 826
rect 225 801 227 804
rect 240 795 242 796
rect 211 792 213 793
rect 240 772 242 775
rect 211 769 213 772
rect 255 762 257 765
rect 63 755 65 759
rect 73 755 75 759
rect 215 756 217 759
rect 407 744 409 747
rect 63 716 65 735
rect 73 716 75 735
rect 104 723 106 726
rect 215 724 217 736
rect 255 730 257 742
rect 328 738 330 741
rect 26 698 28 701
rect 36 698 38 701
rect 215 711 217 714
rect 255 707 257 710
rect 328 706 330 718
rect 407 712 409 724
rect 63 693 65 696
rect 73 693 75 696
rect 104 691 106 703
rect 407 699 409 702
rect 328 693 330 696
rect 422 693 424 694
rect 393 690 395 691
rect 343 687 345 688
rect 314 684 316 685
rect 104 678 106 681
rect 422 670 424 673
rect 393 667 395 670
rect 343 664 345 667
rect 95 661 97 664
rect 105 661 107 664
rect 314 661 316 664
rect 26 639 28 658
rect 36 639 38 658
rect 26 626 28 629
rect 36 626 38 629
rect 437 660 439 663
rect 358 654 360 657
rect 397 654 399 657
rect 318 648 320 651
rect 130 641 132 644
rect 26 618 28 621
rect 36 618 38 621
rect 95 603 97 621
rect 105 603 107 621
rect 130 607 132 621
rect 161 616 163 620
rect 171 616 173 620
rect 318 616 320 628
rect 358 622 360 634
rect 397 622 399 634
rect 437 628 439 640
rect 26 578 28 598
rect 36 578 38 598
rect 130 594 132 597
rect 318 603 320 606
rect 397 609 399 612
rect 437 605 439 608
rect 358 599 360 602
rect 95 590 97 593
rect 105 590 107 593
rect 161 577 163 596
rect 171 577 173 596
rect 95 563 97 566
rect 105 563 107 566
rect 26 554 28 558
rect 36 554 38 558
rect 21 524 23 527
rect 31 524 33 527
rect 326 566 328 569
rect 417 566 419 569
rect 161 554 163 557
rect 171 554 173 557
rect 153 531 155 535
rect 163 531 165 535
rect 326 534 328 546
rect 417 534 419 546
rect 187 531 189 534
rect 95 505 97 523
rect 105 505 107 523
rect 326 521 328 524
rect 417 521 419 524
rect 341 515 343 516
rect 312 512 314 513
rect 95 492 97 495
rect 105 492 107 495
rect 153 492 155 511
rect 163 492 165 511
rect 187 499 189 511
rect 21 465 23 484
rect 31 465 33 484
rect 85 473 87 476
rect 95 473 97 476
rect 21 452 23 455
rect 31 452 33 455
rect 21 444 23 447
rect 31 444 33 447
rect 432 515 434 516
rect 403 512 405 513
rect 341 492 343 495
rect 432 492 434 495
rect 312 489 314 492
rect 403 489 405 492
rect 187 486 189 489
rect 356 482 358 485
rect 447 482 449 485
rect 316 476 318 479
rect 153 469 155 472
rect 163 469 165 472
rect 208 468 210 471
rect 218 468 220 471
rect 120 453 122 456
rect 21 404 23 424
rect 31 404 33 424
rect 85 415 87 433
rect 95 415 97 433
rect 120 419 122 433
rect 158 429 160 433
rect 168 429 170 433
rect 407 476 409 479
rect 243 448 245 451
rect 316 444 318 456
rect 356 450 358 462
rect 316 431 318 434
rect 407 444 409 456
rect 447 450 449 462
rect 407 431 409 434
rect 208 410 210 428
rect 218 410 220 428
rect 243 414 245 428
rect 356 427 358 430
rect 447 427 449 430
rect 120 406 122 409
rect 85 402 87 405
rect 95 402 97 405
rect 158 390 160 409
rect 168 390 170 409
rect 243 401 245 404
rect 331 400 333 403
rect 418 400 420 403
rect 208 397 210 400
rect 218 397 220 400
rect 21 380 23 384
rect 31 380 33 384
rect 76 375 78 378
rect 86 375 88 378
rect 20 351 22 354
rect 30 351 32 354
rect 158 367 160 370
rect 168 367 170 370
rect 331 368 333 380
rect 418 368 420 380
rect 331 355 333 358
rect 418 355 420 358
rect 346 349 348 350
rect 317 346 319 347
rect 197 336 199 340
rect 207 336 209 340
rect 231 336 233 339
rect 76 317 78 335
rect 86 317 88 335
rect 20 292 22 311
rect 30 292 32 311
rect 433 349 435 350
rect 404 346 406 347
rect 346 326 348 329
rect 433 326 435 329
rect 317 323 319 326
rect 404 323 406 326
rect 361 316 363 319
rect 448 316 450 319
rect 76 304 78 307
rect 86 304 88 307
rect 197 297 199 316
rect 207 297 209 316
rect 231 304 233 316
rect 321 310 323 313
rect 83 282 85 285
rect 93 282 95 285
rect 20 279 22 282
rect 30 279 32 282
rect 20 271 22 274
rect 30 271 32 274
rect 20 231 22 251
rect 30 231 32 251
rect 231 291 233 294
rect 408 310 410 313
rect 321 278 323 290
rect 361 284 363 296
rect 197 274 199 277
rect 207 274 209 277
rect 321 265 323 268
rect 118 262 120 265
rect 408 278 410 290
rect 448 284 450 296
rect 408 265 410 268
rect 361 261 363 264
rect 448 261 450 264
rect 203 251 205 254
rect 213 251 215 254
rect 83 224 85 242
rect 93 224 95 242
rect 118 228 120 242
rect 158 237 160 241
rect 168 237 170 241
rect 118 215 120 218
rect 83 211 85 214
rect 93 211 95 214
rect 20 207 22 211
rect 30 207 32 211
rect 158 198 160 217
rect 168 198 170 217
rect 415 237 417 240
rect 238 231 240 234
rect 83 184 85 187
rect 93 184 95 187
rect 22 151 24 154
rect 32 151 34 154
rect 203 193 205 211
rect 213 193 215 211
rect 238 197 240 211
rect 415 205 417 217
rect 333 195 335 198
rect 238 184 240 187
rect 203 180 205 183
rect 213 180 215 183
rect 158 175 160 178
rect 168 175 170 178
rect 415 192 417 195
rect 430 186 432 187
rect 401 183 403 184
rect 333 163 335 175
rect 430 163 432 166
rect 160 152 162 156
rect 170 152 172 156
rect 194 152 196 155
rect 401 160 403 163
rect 445 153 447 156
rect 83 126 85 144
rect 93 126 95 144
rect 333 150 335 153
rect 405 147 407 150
rect 348 144 350 145
rect 319 141 321 142
rect 83 113 85 116
rect 93 113 95 116
rect 160 113 162 132
rect 170 113 172 132
rect 194 120 196 132
rect 348 121 350 124
rect 22 92 24 111
rect 32 92 34 111
rect 77 94 79 97
rect 87 94 89 97
rect 22 79 24 82
rect 32 79 34 82
rect 22 71 24 74
rect 32 71 34 74
rect 319 118 321 121
rect 405 115 407 127
rect 445 121 447 133
rect 363 111 365 114
rect 194 107 196 110
rect 323 105 325 108
rect 219 99 221 102
rect 229 99 231 102
rect 160 90 162 93
rect 170 90 172 93
rect 112 74 114 77
rect 136 73 138 77
rect 146 73 148 77
rect 22 31 24 51
rect 32 31 34 51
rect 77 36 79 54
rect 87 36 89 54
rect 112 40 114 54
rect 405 102 407 105
rect 445 98 447 101
rect 254 79 256 82
rect 323 73 325 85
rect 363 79 365 91
rect 323 60 325 63
rect 136 34 138 53
rect 146 34 148 53
rect 219 41 221 59
rect 229 41 231 59
rect 254 45 256 59
rect 363 56 365 59
rect 112 27 114 30
rect 77 23 79 26
rect 87 23 89 26
rect 254 32 256 35
rect 219 28 221 31
rect 229 28 231 31
rect 136 11 138 14
rect 146 11 148 14
rect 22 7 24 11
rect 32 7 34 11
<< polycontact >>
rect 221 815 225 819
rect 209 793 213 797
rect 238 796 242 800
rect 59 724 63 728
rect 69 717 73 721
rect 211 725 215 729
rect 324 707 328 711
rect 403 713 407 717
rect 100 692 104 696
rect 312 685 316 689
rect 341 688 345 692
rect 391 691 395 695
rect 420 694 424 698
rect 22 640 26 644
rect 32 647 36 651
rect 91 604 95 608
rect 101 610 105 614
rect 126 608 130 612
rect 314 617 318 621
rect 393 623 397 627
rect 22 585 26 589
rect 32 593 36 597
rect 157 585 161 589
rect 167 578 171 582
rect 322 535 326 539
rect 413 535 417 539
rect 91 506 95 510
rect 101 512 105 516
rect 310 513 314 517
rect 339 516 343 520
rect 149 500 153 504
rect 159 493 163 497
rect 183 500 187 504
rect 17 466 21 470
rect 27 473 31 477
rect 401 513 405 517
rect 430 516 434 520
rect 17 411 21 415
rect 27 419 31 423
rect 81 416 85 420
rect 91 422 95 426
rect 116 420 120 424
rect 312 445 316 449
rect 403 445 407 449
rect 204 411 208 415
rect 214 417 218 421
rect 239 415 243 419
rect 154 398 158 402
rect 164 391 168 395
rect 327 369 331 373
rect 414 369 418 373
rect 315 347 319 351
rect 344 350 348 354
rect 72 318 76 322
rect 82 324 86 328
rect 16 293 20 297
rect 26 300 30 304
rect 402 347 406 351
rect 431 350 435 354
rect 193 305 197 309
rect 203 298 207 302
rect 227 305 231 309
rect 16 238 20 242
rect 26 246 30 250
rect 317 279 321 283
rect 404 279 408 283
rect 79 225 83 229
rect 89 231 93 235
rect 114 229 118 233
rect 154 206 158 210
rect 164 199 168 203
rect 199 194 203 198
rect 209 200 213 204
rect 234 198 238 202
rect 411 206 415 210
rect 399 184 403 188
rect 428 187 432 191
rect 329 164 333 168
rect 79 127 83 131
rect 89 133 93 137
rect 317 142 321 146
rect 346 145 350 149
rect 156 121 160 125
rect 166 114 170 118
rect 190 121 194 125
rect 18 93 22 97
rect 28 100 32 104
rect 401 116 405 120
rect 18 38 22 42
rect 28 46 32 50
rect 73 37 77 41
rect 83 43 87 47
rect 108 41 112 45
rect 319 74 323 78
rect 132 42 136 46
rect 142 35 146 39
rect 215 42 219 46
rect 225 48 229 52
rect 250 46 254 50
<< polynpluscontact >>
rect 251 731 255 735
rect 354 623 358 627
rect 433 629 437 633
rect 352 451 356 455
rect 443 451 447 455
rect 357 285 361 289
rect 444 285 448 289
rect 441 122 445 126
rect 359 80 363 84
<< metal1 >>
rect 199 853 253 856
rect 199 777 202 853
rect 220 846 223 853
rect 210 815 221 818
rect 229 818 232 826
rect 229 815 241 818
rect 205 797 208 815
rect 229 814 232 815
rect 220 800 223 804
rect 238 800 241 815
rect 220 797 225 800
rect 205 794 209 797
rect 244 772 247 775
rect 215 769 247 772
rect 58 762 80 765
rect 199 763 215 766
rect 58 755 61 762
rect 77 755 80 762
rect 210 756 213 763
rect 45 724 59 727
rect 68 727 71 735
rect 94 730 104 733
rect 68 724 86 727
rect 45 717 69 720
rect 77 716 80 724
rect 15 704 44 708
rect 21 698 25 704
rect 58 693 61 696
rect 83 695 86 724
rect 99 723 102 730
rect 204 725 211 728
rect 219 728 222 736
rect 244 734 247 769
rect 250 762 253 853
rect 381 751 435 754
rect 244 731 251 734
rect 259 734 262 742
rect 302 745 356 748
rect 259 731 278 734
rect 259 730 262 731
rect 219 725 234 728
rect 219 724 222 725
rect 210 707 213 714
rect 250 707 253 710
rect 210 704 225 707
rect 108 696 111 703
rect 230 704 253 707
rect 57 690 62 693
rect 79 692 100 695
rect 108 693 148 696
rect 6 647 32 651
rect 6 623 9 647
rect 39 644 43 658
rect 6 589 9 618
rect 12 640 22 644
rect 30 640 70 644
rect 30 639 34 640
rect 12 597 15 635
rect 21 625 25 629
rect 39 625 43 629
rect 21 622 43 625
rect 21 618 25 622
rect 66 607 70 640
rect 83 614 86 692
rect 108 691 111 693
rect 99 677 102 681
rect 99 674 109 677
rect 90 668 123 671
rect 302 669 305 745
rect 323 738 326 745
rect 313 707 324 710
rect 332 710 335 718
rect 332 707 344 710
rect 308 689 311 707
rect 332 706 335 707
rect 323 692 326 696
rect 341 692 344 707
rect 323 689 328 692
rect 308 686 312 689
rect 90 661 93 668
rect 120 651 123 668
rect 347 664 350 667
rect 318 661 350 664
rect 302 655 318 658
rect 120 648 128 651
rect 125 641 128 648
rect 313 648 316 655
rect 83 611 101 614
rect 109 612 112 621
rect 134 612 137 621
rect 156 623 178 626
rect 156 616 159 623
rect 175 616 178 623
rect 307 617 314 620
rect 322 620 325 628
rect 347 626 350 661
rect 353 654 356 745
rect 381 675 384 751
rect 402 744 405 751
rect 387 713 403 716
rect 411 716 414 724
rect 411 713 423 716
rect 387 704 390 713
rect 411 712 414 713
rect 387 695 390 699
rect 402 698 405 702
rect 420 698 423 713
rect 402 695 407 698
rect 387 692 391 695
rect 426 670 429 673
rect 397 667 429 670
rect 381 661 397 664
rect 392 654 395 661
rect 347 623 354 626
rect 362 626 365 634
rect 362 623 381 626
rect 362 622 365 623
rect 322 617 337 620
rect 386 623 393 626
rect 401 626 404 634
rect 426 632 429 667
rect 432 660 435 751
rect 426 629 433 632
rect 441 632 444 640
rect 441 629 450 632
rect 441 628 444 629
rect 401 623 416 626
rect 401 622 404 623
rect 322 616 325 617
rect 109 609 126 612
rect 66 604 76 607
rect 81 604 91 607
rect 109 607 112 609
rect 134 609 143 612
rect 134 607 137 609
rect 100 604 112 607
rect 100 603 103 604
rect 12 593 32 597
rect 39 589 43 598
rect 6 585 22 589
rect 30 585 65 589
rect 30 578 34 585
rect 61 581 65 585
rect 90 587 93 593
rect 109 587 112 593
rect 125 587 128 597
rect 90 584 128 587
rect 140 588 143 609
rect 313 599 316 606
rect 392 605 395 612
rect 432 605 435 608
rect 392 602 407 605
rect 353 599 356 602
rect 412 602 435 605
rect 313 596 328 599
rect 140 585 157 588
rect 166 588 169 596
rect 333 596 356 599
rect 166 585 187 588
rect 58 578 167 581
rect 175 577 178 585
rect 88 572 94 575
rect 300 573 354 576
rect 90 563 93 572
rect 21 550 25 558
rect 39 552 43 558
rect 156 554 159 557
rect 39 550 44 552
rect 21 547 44 550
rect 155 551 160 554
rect 148 538 185 541
rect 10 530 39 534
rect 148 531 151 538
rect 167 531 170 538
rect 16 524 20 530
rect 182 531 185 538
rect 82 513 101 516
rect 109 514 112 523
rect 109 511 120 514
rect 46 506 62 509
rect 67 506 91 509
rect 109 509 112 511
rect 100 506 112 509
rect 1 473 27 477
rect 1 450 4 473
rect 34 470 38 484
rect 46 470 49 506
rect 1 415 4 445
rect 12 466 17 470
rect 25 466 49 470
rect 25 465 29 466
rect 7 423 10 465
rect 16 451 20 455
rect 34 451 38 455
rect 16 448 38 451
rect 16 444 20 448
rect 7 419 27 423
rect 34 415 38 424
rect 73 426 76 506
rect 100 505 103 506
rect 90 489 93 495
rect 109 489 112 495
rect 117 496 120 511
rect 138 500 149 503
rect 158 503 161 511
rect 191 504 194 511
rect 158 500 183 503
rect 191 501 200 504
rect 117 493 159 496
rect 167 492 170 500
rect 191 499 194 501
rect 90 486 112 489
rect 80 480 113 483
rect 80 473 83 480
rect 110 463 113 480
rect 148 469 151 472
rect 182 469 185 489
rect 147 466 185 469
rect 110 460 118 463
rect 115 453 118 460
rect 73 423 91 426
rect 99 424 102 433
rect 124 424 127 433
rect 153 436 175 439
rect 153 429 156 436
rect 172 429 175 436
rect 99 421 116 424
rect 60 416 81 419
rect 99 419 102 421
rect 124 421 133 424
rect 197 421 200 501
rect 300 497 303 573
rect 321 566 324 573
rect 311 535 322 538
rect 330 538 333 546
rect 330 535 342 538
rect 306 517 309 535
rect 330 534 333 535
rect 321 520 324 524
rect 339 520 342 535
rect 321 517 326 520
rect 306 514 310 517
rect 345 492 348 495
rect 316 489 348 492
rect 300 483 316 486
rect 203 475 236 478
rect 203 468 206 475
rect 233 458 236 475
rect 311 476 314 483
rect 233 455 241 458
rect 238 448 241 455
rect 305 445 312 448
rect 320 448 323 456
rect 345 454 348 489
rect 351 482 354 573
rect 391 573 445 576
rect 391 497 394 573
rect 412 566 415 573
rect 402 535 413 538
rect 421 538 424 546
rect 421 535 433 538
rect 397 517 400 535
rect 421 534 424 535
rect 412 520 415 524
rect 430 520 433 535
rect 412 517 417 520
rect 397 514 401 517
rect 436 492 439 495
rect 407 489 439 492
rect 391 483 407 486
rect 402 476 405 483
rect 345 451 352 454
rect 360 454 363 462
rect 360 451 369 454
rect 360 450 363 451
rect 320 445 335 448
rect 366 448 369 451
rect 366 445 391 448
rect 320 444 323 445
rect 396 445 403 448
rect 411 448 414 456
rect 436 454 439 489
rect 442 482 445 573
rect 436 451 443 454
rect 451 454 454 462
rect 451 451 460 454
rect 451 450 454 451
rect 411 445 426 448
rect 411 444 414 445
rect 124 419 127 421
rect 90 416 102 419
rect 90 415 93 416
rect 1 411 17 415
rect 25 411 50 415
rect 25 404 29 411
rect 47 393 50 411
rect 80 399 83 405
rect 99 399 102 405
rect 115 399 118 409
rect 80 396 118 399
rect 130 401 133 421
rect 196 418 214 421
rect 222 419 225 428
rect 247 419 250 428
rect 311 427 314 434
rect 351 427 354 430
rect 311 424 326 427
rect 331 424 354 427
rect 402 427 405 434
rect 442 427 445 430
rect 402 424 417 427
rect 422 424 445 427
rect 222 416 239 419
rect 130 398 154 401
rect 163 401 166 409
rect 192 411 204 414
rect 222 414 225 416
rect 247 416 256 419
rect 247 414 250 416
rect 213 411 225 414
rect 192 401 195 411
rect 213 410 216 411
rect 305 407 359 410
rect 163 398 195 401
rect 47 390 71 393
rect 146 393 164 394
rect 76 391 164 393
rect 76 390 149 391
rect 172 390 175 398
rect 203 394 206 400
rect 222 394 225 400
rect 238 394 241 404
rect 203 391 241 394
rect 16 376 20 384
rect 69 384 75 387
rect 34 378 38 384
rect 34 376 39 378
rect 16 373 39 376
rect 71 375 74 384
rect 153 367 156 370
rect 152 364 157 367
rect 9 357 38 361
rect 15 351 19 357
rect 192 343 229 346
rect 63 325 82 328
rect 90 326 93 335
rect 192 336 195 343
rect 211 336 214 343
rect 226 336 229 343
rect 305 331 308 407
rect 326 400 329 407
rect 316 369 327 372
rect 335 372 338 380
rect 335 369 347 372
rect 311 351 314 369
rect 335 368 338 369
rect 326 354 329 358
rect 344 354 347 369
rect 326 351 331 354
rect 311 348 315 351
rect 350 326 353 329
rect 90 323 143 326
rect 321 323 353 326
rect 46 318 72 321
rect 90 321 93 323
rect 81 318 93 321
rect 0 300 26 304
rect 0 284 3 300
rect 33 297 37 311
rect 46 297 50 318
rect 0 242 3 279
rect 11 293 16 297
rect 24 293 50 297
rect 24 292 28 293
rect 6 250 9 292
rect 15 278 19 282
rect 33 278 37 282
rect 15 275 37 278
rect 15 271 19 275
rect 6 246 26 250
rect 33 242 37 251
rect 0 238 16 242
rect 24 238 47 242
rect 24 231 28 238
rect 59 228 62 318
rect 81 317 84 318
rect 71 301 74 307
rect 90 301 93 307
rect 71 298 93 301
rect 140 301 143 323
rect 305 317 321 320
rect 184 305 193 308
rect 202 308 205 316
rect 235 309 238 316
rect 316 310 319 317
rect 202 305 227 308
rect 235 306 244 309
rect 140 298 203 301
rect 211 297 214 305
rect 235 304 238 306
rect 78 289 111 292
rect 78 282 81 289
rect 108 272 111 289
rect 192 274 195 277
rect 226 274 229 294
rect 108 269 116 272
rect 191 271 229 274
rect 113 262 116 269
rect 241 268 244 306
rect 310 279 317 282
rect 325 282 328 290
rect 350 288 353 323
rect 356 316 359 407
rect 392 407 446 410
rect 392 331 395 407
rect 413 400 416 407
rect 403 369 414 372
rect 422 372 425 380
rect 422 369 434 372
rect 398 351 401 369
rect 422 368 425 369
rect 413 354 416 358
rect 431 354 434 369
rect 413 351 418 354
rect 398 348 402 351
rect 437 326 440 329
rect 408 323 440 326
rect 392 317 408 320
rect 403 310 406 317
rect 350 285 357 288
rect 365 288 368 296
rect 365 285 387 288
rect 365 284 368 285
rect 325 279 340 282
rect 384 282 387 285
rect 384 279 392 282
rect 325 278 328 279
rect 397 279 404 282
rect 412 282 415 290
rect 437 288 440 323
rect 443 316 446 407
rect 437 285 444 288
rect 452 288 455 296
rect 452 285 461 288
rect 452 284 455 285
rect 412 279 427 282
rect 412 278 415 279
rect 192 265 244 268
rect 70 232 89 235
rect 97 233 100 242
rect 122 233 125 242
rect 153 244 175 247
rect 153 237 156 244
rect 172 237 175 244
rect 97 230 114 233
rect 59 225 79 228
rect 97 228 100 230
rect 122 230 131 233
rect 122 228 125 230
rect 88 225 100 228
rect 15 203 19 211
rect 33 205 37 211
rect 33 203 38 205
rect 15 200 38 203
rect 11 157 40 161
rect 17 151 21 157
rect 59 137 62 225
rect 88 224 91 225
rect 78 208 81 214
rect 97 208 100 214
rect 113 208 116 218
rect 78 205 116 208
rect 128 209 131 230
rect 128 206 154 209
rect 163 209 166 217
rect 163 206 181 209
rect 71 199 164 202
rect 172 198 175 206
rect 76 193 82 196
rect 178 197 181 206
rect 192 204 195 265
rect 316 261 319 268
rect 356 261 359 264
rect 198 258 231 261
rect 316 258 331 261
rect 198 251 201 258
rect 228 241 231 258
rect 336 258 359 261
rect 403 261 406 268
rect 443 261 446 264
rect 403 258 418 261
rect 423 258 446 261
rect 389 244 443 247
rect 228 238 236 241
rect 233 231 236 238
rect 192 201 209 204
rect 217 202 220 211
rect 242 202 245 211
rect 217 199 234 202
rect 178 194 199 197
rect 217 197 220 199
rect 242 199 249 202
rect 307 202 361 205
rect 242 197 245 199
rect 208 194 220 197
rect 208 193 211 194
rect 78 184 81 193
rect 153 175 156 178
rect 198 177 201 183
rect 217 177 220 183
rect 233 177 236 187
rect 152 172 157 175
rect 198 174 236 177
rect 155 159 192 162
rect 155 152 158 159
rect 174 152 177 159
rect 189 152 192 159
rect 59 134 89 137
rect 97 135 100 144
rect 97 132 132 135
rect 59 127 79 130
rect 97 130 100 132
rect 88 127 100 130
rect 2 100 28 104
rect 2 79 5 100
rect 35 97 39 111
rect 59 97 62 127
rect 88 126 91 127
rect 78 110 81 116
rect 97 110 100 116
rect 129 117 132 132
rect 148 121 156 124
rect 165 124 168 132
rect 198 125 201 132
rect 307 126 310 202
rect 328 195 331 202
rect 318 164 329 167
rect 337 167 340 175
rect 337 164 349 167
rect 337 163 340 164
rect 313 146 316 162
rect 328 149 331 153
rect 346 149 349 164
rect 328 146 333 149
rect 313 143 317 146
rect 165 121 190 124
rect 198 122 207 125
rect 129 114 166 117
rect 174 113 177 121
rect 198 120 201 122
rect 78 107 100 110
rect 2 42 5 74
rect 13 93 18 97
rect 26 93 62 97
rect 26 92 30 93
rect 8 50 11 92
rect 17 78 21 82
rect 35 78 39 82
rect 17 75 39 78
rect 17 71 21 75
rect 59 63 62 93
rect 72 101 105 104
rect 72 94 75 101
rect 102 84 105 101
rect 155 90 158 93
rect 189 90 192 110
rect 154 87 192 90
rect 102 81 110 84
rect 107 74 110 81
rect 131 80 153 83
rect 131 73 134 80
rect 150 73 153 80
rect 51 60 62 63
rect 8 46 28 50
rect 35 42 39 51
rect 2 38 18 42
rect 26 38 45 42
rect 26 31 30 38
rect 17 3 21 11
rect 35 5 39 11
rect 42 11 45 38
rect 51 40 54 60
rect 63 44 83 47
rect 91 45 94 54
rect 116 45 119 54
rect 91 42 108 45
rect 51 37 73 40
rect 91 40 94 42
rect 116 42 132 45
rect 141 45 144 53
rect 204 52 207 122
rect 352 121 355 124
rect 323 118 355 121
rect 307 112 323 115
rect 214 106 247 109
rect 214 99 217 106
rect 244 89 247 106
rect 318 105 321 112
rect 244 86 252 89
rect 249 79 252 86
rect 312 74 319 77
rect 327 77 330 85
rect 352 83 355 118
rect 358 111 361 202
rect 389 168 392 244
rect 410 237 413 244
rect 395 206 411 209
rect 419 209 422 217
rect 419 206 431 209
rect 395 203 398 206
rect 419 205 422 206
rect 395 188 398 198
rect 410 191 413 195
rect 428 191 431 206
rect 410 188 415 191
rect 395 185 399 188
rect 434 163 437 166
rect 405 160 437 163
rect 389 154 405 157
rect 400 147 403 154
rect 394 116 401 119
rect 409 119 412 127
rect 434 125 437 160
rect 440 153 443 244
rect 434 122 441 125
rect 449 125 452 133
rect 449 122 458 125
rect 449 121 452 122
rect 409 116 424 119
rect 409 115 412 116
rect 352 80 359 83
rect 367 83 370 91
rect 389 83 392 114
rect 400 98 403 105
rect 440 98 443 101
rect 400 95 415 98
rect 420 95 443 98
rect 367 80 392 83
rect 367 79 370 80
rect 327 74 342 77
rect 327 73 330 74
rect 204 49 225 52
rect 233 50 236 59
rect 258 50 261 59
rect 318 56 321 63
rect 358 56 361 59
rect 318 53 333 56
rect 338 53 361 56
rect 233 47 250 50
rect 141 42 215 45
rect 233 45 236 47
rect 258 47 267 50
rect 258 45 261 47
rect 224 42 236 45
rect 116 40 119 42
rect 82 37 94 40
rect 82 36 85 37
rect 122 35 142 38
rect 72 20 75 26
rect 91 20 94 26
rect 107 20 110 30
rect 72 17 110 20
rect 122 11 125 35
rect 150 34 153 42
rect 224 41 227 42
rect 214 25 217 31
rect 233 25 236 31
rect 249 25 252 35
rect 214 22 252 25
rect 131 11 134 14
rect 42 8 125 11
rect 130 8 135 11
rect 35 3 40 5
rect 17 0 40 3
<< m2contact >>
rect 225 795 230 800
rect 44 704 49 709
rect 234 725 239 730
rect 225 702 230 707
rect 148 693 153 698
rect 328 687 333 692
rect 387 699 392 704
rect 407 693 412 698
rect 337 617 342 622
rect 381 621 386 626
rect 416 623 421 628
rect 76 602 81 607
rect 407 600 412 605
rect 328 594 333 599
rect 187 585 192 590
rect 53 576 58 581
rect 44 547 49 552
rect 39 530 44 535
rect 77 513 82 518
rect 62 506 67 511
rect 55 416 60 421
rect 326 515 331 520
rect 397 535 402 540
rect 417 515 422 520
rect 335 445 340 450
rect 391 443 396 448
rect 426 445 431 450
rect 326 422 331 427
rect 417 422 422 427
rect 256 416 261 421
rect 71 390 76 395
rect 39 373 44 378
rect 38 357 43 362
rect 58 325 63 330
rect 331 349 336 354
rect 47 238 52 243
rect 179 305 184 310
rect 398 369 403 374
rect 418 349 423 354
rect 340 279 345 284
rect 392 277 397 282
rect 427 279 432 284
rect 65 232 70 237
rect 38 200 43 205
rect 40 157 45 162
rect 65 199 71 205
rect 331 256 336 261
rect 418 256 423 261
rect 143 121 148 126
rect 333 144 338 149
rect 58 44 63 49
rect 415 186 420 191
rect 389 114 394 119
rect 424 116 429 121
rect 415 93 420 98
rect 342 74 347 79
rect 333 51 338 56
rect 40 0 45 5
<< psm12contact >>
rect 133 500 138 505
<< ndm12contact >>
rect 205 772 210 777
rect 234 775 239 780
rect 308 664 313 669
rect 337 667 342 672
rect 387 670 392 675
rect 416 673 421 678
rect 306 492 311 497
rect 335 495 340 500
rect 397 492 402 497
rect 426 495 431 500
rect 311 326 316 331
rect 340 329 345 334
rect 398 326 403 331
rect 427 329 432 334
rect 313 121 318 126
rect 342 124 347 129
rect 395 163 400 168
rect 424 166 429 171
<< metal2 >>
rect 199 772 205 777
rect 199 728 202 772
rect 227 707 230 795
rect 234 730 237 775
rect 46 552 49 704
rect 278 699 387 702
rect 278 696 281 699
rect 153 693 281 696
rect 41 378 44 530
rect 55 421 58 576
rect 78 518 81 602
rect 148 515 151 693
rect 302 664 308 669
rect 302 620 305 664
rect 330 599 333 687
rect 381 670 387 675
rect 337 622 340 667
rect 381 626 384 670
rect 409 605 412 693
rect 416 628 419 673
rect 133 512 151 515
rect 189 563 192 585
rect 189 560 400 563
rect 40 205 43 357
rect 64 335 67 506
rect 133 505 136 512
rect 58 332 67 335
rect 58 330 64 332
rect 73 240 76 390
rect 189 317 192 560
rect 397 540 400 560
rect 300 492 306 497
rect 300 448 303 492
rect 328 427 331 515
rect 335 450 338 495
rect 391 492 397 497
rect 391 448 394 492
rect 419 427 422 515
rect 426 450 429 495
rect 181 314 192 317
rect 258 387 261 416
rect 258 384 401 387
rect 181 310 184 314
rect 49 202 52 238
rect 65 237 76 240
rect 49 199 65 202
rect 42 5 45 157
rect 65 59 68 199
rect 258 168 261 384
rect 398 374 401 384
rect 305 326 311 331
rect 305 282 308 326
rect 333 261 336 349
rect 340 284 343 329
rect 392 326 398 331
rect 392 282 395 326
rect 420 261 423 349
rect 427 284 430 329
rect 143 165 261 168
rect 143 126 146 165
rect 389 163 395 168
rect 307 121 313 126
rect 307 77 310 121
rect 60 56 68 59
rect 335 56 338 144
rect 342 79 345 124
rect 389 119 392 163
rect 417 98 420 186
rect 424 121 427 166
rect 60 49 63 56
<< m123contact >>
rect 205 815 210 820
rect 40 724 45 729
rect 199 723 204 728
rect 40 715 45 720
rect 308 707 313 712
rect 12 635 17 640
rect 4 618 9 623
rect 7 465 12 470
rect -1 445 4 450
rect 302 615 307 620
rect 6 292 11 297
rect -2 279 3 284
rect 306 535 311 540
rect 300 443 305 448
rect 249 199 254 204
rect 8 92 13 97
rect 0 74 5 79
rect 311 369 316 374
rect 305 277 310 282
rect 395 198 400 203
rect 313 162 318 167
rect 307 72 312 77
<< metal3 >>
rect 191 815 205 820
rect 191 729 195 815
rect 45 724 195 729
rect 199 720 204 723
rect 45 715 204 720
rect 294 707 308 711
rect 294 640 298 707
rect 17 636 298 640
rect 9 619 298 622
rect 9 618 302 619
rect 294 615 302 618
rect 286 535 306 538
rect 286 470 289 535
rect 12 467 289 470
rect 4 445 300 448
rect 290 370 311 373
rect 290 297 293 370
rect 11 294 293 297
rect 3 279 305 282
rect 254 199 395 202
rect 297 162 313 165
rect 297 97 300 162
rect 13 94 300 97
rect 5 74 307 77
<< labels >>
rlabel metal1 98 732 98 732 4 vdd
rlabel metal1 105 675 105 675 1 gnd
rlabel metal1 114 694 114 694 7 c1
rlabel metal1 100 585 100 585 1 gnd
rlabel metal1 105 669 105 669 5 vdd
rlabel metal1 80 693 80 693 3 g0_bar
rlabel metal1 67 605 67 605 3 p1_bar
rlabel metal1 167 624 167 624 5 vdd
rlabel metal1 158 552 158 552 1 gnd
rlabel metal1 67 579 67 579 3 g1_bar
rlabel metal1 181 587 181 587 7 c2
rlabel metal1 91 574 91 574 5 vdd
rlabel metal1 100 487 100 487 1 gnd
rlabel metal1 54 507 54 507 3 p2_bar
rlabel metal1 90 397 90 397 1 gnd
rlabel metal1 95 481 95 481 5 vdd
rlabel metal1 163 540 163 540 1 vdd
rlabel metal1 168 467 168 467 1 gnd
rlabel metal1 155 365 155 365 1 gnd
rlabel metal1 164 437 164 437 5 vdd
rlabel metal1 218 477 218 477 1 vdd
rlabel metal1 219 392 219 392 1 gnd
rlabel metal1 71 385 71 385 1 vdd
rlabel metal1 80 299 80 299 1 gnd
rlabel metal1 91 290 91 290 1 vdd
rlabel metal1 96 206 96 206 1 gnd
rlabel metal1 163 245 163 245 1 vdd
rlabel metal1 155 173 155 173 1 gnd
rlabel metal1 253 417 253 417 7 c3
rlabel metal1 207 345 207 345 1 vdd
rlabel metal1 212 273 212 273 1 gnd
rlabel metal1 217 175 217 175 1 gnd
rlabel metal1 215 259 215 259 1 vdd
rlabel metal1 249 200 249 200 1 c4
rlabel metal1 80 200 80 200 1 g3_bar
rlabel metal1 78 194 78 194 1 vdd
rlabel metal1 86 108 86 108 1 gnd
rlabel metal1 60 128 60 128 1 p4_bar
rlabel metal1 87 102 87 102 1 vdd
rlabel metal1 92 18 92 18 1 gnd
rlabel metal1 50 9 50 9 1 g4_bar
rlabel metal1 171 160 171 160 1 vdd
rlabel metal1 173 88 173 88 1 gnd
rlabel metal1 131 9 131 9 1 gnd
rlabel metal1 142 81 142 81 1 vdd
rlabel metal1 234 23 234 23 1 gnd
rlabel metal1 230 107 230 107 1 vdd
rlabel metal1 264 48 264 48 7 c5
rlabel metal1 31 706 31 706 5 vdd
rlabel metal1 32 624 32 624 1 gnd
rlabel metal1 13 617 13 617 1 b1
rlabel metal1 7 617 7 617 3 a1
rlabel metal1 69 763 69 763 5 vdd
rlabel metal1 59 691 59 691 1 gnd
rlabel metal1 53 725 53 725 1 a0
rlabel metal1 53 718 53 718 1 b0
rlabel metal1 50 391 50 391 1 g2_bar
rlabel metal1 26 532 26 532 1 vdd
rlabel metal1 27 449 27 449 1 gnd
rlabel metal1 8 441 8 441 1 b2
rlabel metal1 2 441 2 441 3 a2
rlabel metal1 55 319 55 319 1 p3_bar
rlabel metal1 24 359 24 359 1 vdd
rlabel metal1 26 276 26 276 1 gnd
rlabel metal1 8 274 8 274 1 b3
rlabel metal1 1 274 1 274 3 a3
rlabel metal1 24 158 24 158 1 vdd
rlabel metal1 28 76 28 76 1 gnd
rlabel metal1 9 72 9 72 1 b4
rlabel metal1 3 72 3 72 3 a4
rlabel metal1 237 706 237 706 1 gnd
rlabel metal1 221 855 221 855 5 vdd
rlabel metal1 271 732 271 732 1 s0
rlabel metal1 324 746 324 746 1 vdd
rlabel metal1 335 597 335 597 1 gnd
rlabel metal1 372 624 372 624 7 p1
rlabel metal1 447 630 447 630 7 s1
rlabel metal1 415 603 415 603 1 gnd
rlabel metal1 404 753 404 753 1 vdd
rlabel metal1 322 575 322 575 1 vdd
rlabel metal1 337 425 337 425 1 gnd
rlabel metal1 367 452 367 452 1 p2
rlabel metal1 428 425 428 425 1 gnd
rlabel metal1 416 575 416 575 1 vdd
rlabel metal1 330 408 330 408 1 vdd
rlabel metal1 325 259 325 259 1 gnd
rlabel metal1 372 286 372 286 1 p3
rlabel metal1 414 260 414 260 1 gnd
rlabel metal1 415 408 415 408 1 vdd
rlabel metal1 458 287 458 287 7 s3
rlabel metal1 333 204 333 204 1 vdd
rlabel metal1 341 54 341 54 1 gnd
rlabel metal1 373 81 373 81 1 p4
rlabel metal1 412 245 412 245 1 vdd
rlabel metal1 426 96 426 96 1 gnd
rlabel metal1 454 123 454 123 1 s4
rlabel metal1 457 452 457 452 7 s2
rlabel metal1 205 765 205 765 1 vdd
rlabel metal1 308 657 308 657 1 vdd
rlabel metal1 387 663 387 663 1 vdd
rlabel metal1 307 484 307 484 1 vdd
rlabel metal1 397 484 397 484 1 vdd
rlabel metal1 311 319 311 319 1 vdd
rlabel metal1 398 319 398 319 1 vdd
rlabel metal1 312 114 312 114 1 vdd
rlabel metal1 395 155 395 155 1 vdd
<< end >>
