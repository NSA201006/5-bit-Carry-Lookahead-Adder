magic
tech scmos
timestamp 1764648271
<< nwell >>
rect 15 118 39 150
rect 92 118 116 150
rect 5 28 29 60
rect 45 34 69 66
rect 82 28 106 60
rect 122 34 146 66
<< ntransistor >>
rect 26 102 28 112
rect 103 102 105 112
rect 12 70 14 90
rect 41 73 43 93
rect 89 70 91 90
rect 118 73 120 93
rect 16 12 18 22
rect 56 8 58 28
rect 93 12 95 22
rect 133 8 135 28
<< ptransistor >>
rect 26 124 28 144
rect 103 124 105 144
rect 16 34 18 54
rect 56 40 58 60
rect 93 34 95 54
rect 133 40 135 60
<< ndiffusion >>
rect 21 106 26 112
rect 25 102 26 106
rect 28 108 29 112
rect 28 102 33 108
rect 98 106 103 112
rect 102 102 103 106
rect 105 108 106 112
rect 105 102 110 108
rect 6 75 12 90
rect 11 70 12 75
rect 14 74 19 90
rect 14 70 15 74
rect 35 78 41 93
rect 40 73 41 78
rect 43 77 48 93
rect 43 73 44 77
rect 83 75 89 90
rect 88 70 89 75
rect 91 74 96 90
rect 91 70 92 74
rect 112 78 118 93
rect 117 73 118 78
rect 120 77 125 93
rect 120 73 121 77
rect 11 16 16 22
rect 15 12 16 16
rect 18 18 19 22
rect 18 12 23 18
rect 51 12 56 28
rect 55 8 56 12
rect 58 24 59 28
rect 58 8 63 24
rect 88 16 93 22
rect 92 12 93 16
rect 95 18 96 22
rect 95 12 100 18
rect 128 12 133 28
rect 132 8 133 12
rect 135 24 136 28
rect 135 8 140 24
<< pdiffusion >>
rect 25 140 26 144
rect 21 124 26 140
rect 28 128 33 144
rect 28 124 29 128
rect 102 140 103 144
rect 98 124 103 140
rect 105 128 110 144
rect 105 124 106 128
rect 55 56 56 60
rect 15 50 16 54
rect 11 34 16 50
rect 18 38 23 54
rect 51 40 56 56
rect 58 44 63 60
rect 132 56 133 60
rect 58 40 59 44
rect 92 50 93 54
rect 18 34 19 38
rect 88 34 93 50
rect 95 38 100 54
rect 128 40 133 56
rect 135 44 140 60
rect 135 40 136 44
rect 95 34 96 38
<< ndcontact >>
rect 21 102 25 106
rect 29 108 33 112
rect 98 102 102 106
rect 106 108 110 112
rect 15 70 19 74
rect 44 73 48 77
rect 92 70 96 74
rect 121 73 125 77
rect 11 12 15 16
rect 19 18 23 22
rect 51 8 55 12
rect 59 24 63 28
rect 88 12 92 16
rect 96 18 100 22
rect 128 8 132 12
rect 136 24 140 28
<< pdcontact >>
rect 21 140 25 144
rect 29 124 33 128
rect 98 140 102 144
rect 106 124 110 128
rect 51 56 55 60
rect 11 50 15 54
rect 128 56 132 60
rect 59 40 63 44
rect 88 50 92 54
rect 19 34 23 38
rect 136 40 140 44
rect 96 34 100 38
<< polysilicon >>
rect 26 144 28 147
rect 103 144 105 147
rect 26 112 28 124
rect 103 112 105 124
rect 26 99 28 102
rect 103 99 105 102
rect 41 93 43 94
rect 12 90 14 91
rect 118 93 120 94
rect 89 90 91 91
rect 41 70 43 73
rect 118 70 120 73
rect 12 67 14 70
rect 89 67 91 70
rect 56 60 58 63
rect 133 60 135 63
rect 16 54 18 57
rect 93 54 95 57
rect 16 22 18 34
rect 56 28 58 40
rect 16 9 18 12
rect 93 22 95 34
rect 133 28 135 40
rect 93 9 95 12
rect 56 5 58 8
rect 133 5 135 8
<< polycontact >>
rect 22 113 26 117
rect 99 113 103 117
rect 10 91 14 95
rect 39 94 43 98
rect 87 91 91 95
rect 116 94 120 98
rect 12 23 16 27
rect 89 23 93 27
<< polynpluscontact >>
rect 52 29 56 33
rect 129 29 133 33
<< metal1 >>
rect 0 151 131 154
rect 0 64 3 151
rect 21 144 24 151
rect 6 113 22 116
rect 30 116 33 124
rect 30 113 42 116
rect 6 95 9 113
rect 30 112 33 113
rect 21 98 24 102
rect 39 98 42 113
rect 21 95 26 98
rect 6 92 10 95
rect 45 70 48 73
rect 16 67 48 70
rect 0 61 16 64
rect 11 54 14 61
rect 5 23 12 26
rect 20 26 23 34
rect 45 32 48 67
rect 51 60 54 151
rect 77 64 80 151
rect 98 144 101 151
rect 83 113 99 116
rect 107 116 110 124
rect 107 113 119 116
rect 83 95 86 113
rect 107 112 110 113
rect 98 98 101 102
rect 116 98 119 113
rect 98 95 103 98
rect 83 92 87 95
rect 122 70 125 73
rect 93 67 125 70
rect 77 61 93 64
rect 88 54 91 61
rect 45 29 52 32
rect 60 32 63 40
rect 60 29 73 32
rect 60 28 63 29
rect 20 23 35 26
rect 70 26 73 29
rect 70 23 77 26
rect 20 22 23 23
rect 82 23 89 26
rect 97 26 100 34
rect 122 32 125 67
rect 128 60 131 151
rect 122 29 129 32
rect 137 32 140 40
rect 137 29 146 32
rect 137 28 140 29
rect 97 23 112 26
rect 97 22 100 23
rect 11 5 14 12
rect 51 5 54 8
rect 88 5 91 12
rect 128 5 131 8
rect 11 2 26 5
rect 31 2 103 5
rect 108 2 131 5
<< m2contact >>
rect 26 93 31 98
rect 0 21 5 26
rect 103 93 108 98
rect 35 23 40 28
rect 77 21 82 26
rect 112 23 117 28
rect 26 0 31 5
rect 103 0 108 5
<< ndm12contact >>
rect 6 70 11 75
rect 35 73 40 78
rect 83 70 88 75
rect 112 73 117 78
<< metal2 >>
rect 0 70 6 75
rect 0 26 3 70
rect 28 5 31 93
rect 35 28 38 73
rect 77 70 83 75
rect 77 26 80 70
rect 105 5 108 93
rect 112 28 115 73
<< labels >>
rlabel metal1 66 152 66 152 5 vdd
rlabel metal1 73 3 73 3 1 gnd
rlabel metal1 7 24 7 24 1 A
rlabel metal1 8 115 8 115 1 B
rlabel metal1 85 114 85 114 1 C
rlabel metal1 143 30 143 30 7 S
<< end >>
